magic
tech sky130A
magscale 1 2
timestamp 1745668590
<< nwell >>
rect 1066 2159 18898 17425
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 842 2128 18860 17456
<< obsm2 >>
rect 846 2139 18564 17445
<< metal3 >>
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 0 12248 800 12368
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 0 6808 800 6928
rect 0 6128 800 6248
rect 0 5448 800 5568
rect 0 4768 800 4888
<< obsm3 >>
rect 798 15168 17458 17441
rect 880 14888 17458 15168
rect 798 14488 17458 14888
rect 880 14208 17458 14488
rect 798 13808 17458 14208
rect 880 13528 17458 13808
rect 798 13128 17458 13528
rect 880 12848 17458 13128
rect 798 12448 17458 12848
rect 880 12168 17458 12448
rect 798 11768 17458 12168
rect 880 11488 17458 11768
rect 798 11088 17458 11488
rect 880 10808 17458 11088
rect 798 10408 17458 10808
rect 880 10128 17458 10408
rect 798 9728 17458 10128
rect 880 9448 17458 9728
rect 798 9048 17458 9448
rect 880 8768 17458 9048
rect 798 8368 17458 8768
rect 880 8088 17458 8368
rect 798 7688 17458 8088
rect 880 7408 17458 7688
rect 798 7008 17458 7408
rect 880 6728 17458 7008
rect 798 6328 17458 6728
rect 880 6048 17458 6328
rect 798 5648 17458 6048
rect 880 5368 17458 5648
rect 798 4968 17458 5368
rect 880 4688 17458 4968
rect 798 2143 17458 4688
<< metal4 >>
rect 3163 2128 3483 17456
rect 3823 2128 4143 17456
rect 7602 2128 7922 17456
rect 8262 2128 8582 17456
rect 12041 2128 12361 17456
rect 12701 2128 13021 17456
rect 16480 2128 16800 17456
rect 17140 2128 17460 17456
<< metal5 >>
rect 1056 16004 18908 16324
rect 1056 15344 18908 15664
rect 1056 12196 18908 12516
rect 1056 11536 18908 11856
rect 1056 8388 18908 8708
rect 1056 7728 18908 8048
rect 1056 4580 18908 4900
rect 1056 3920 18908 4240
<< labels >>
rlabel metal4 s 3823 2128 4143 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8262 2128 8582 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12701 2128 13021 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17140 2128 17460 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4580 18908 4900 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8388 18908 8708 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12196 18908 12516 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16004 18908 16324 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3163 2128 3483 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3920 18908 4240 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7728 18908 8048 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11536 18908 11856 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15344 18908 15664 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 4768 800 4888 6 x[0]
port 3 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 x[1]
port 4 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 x[2]
port 5 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 x[3]
port 6 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 x[4]
port 7 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 x[5]
port 8 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 x[6]
port 9 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 x[7]
port 10 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 y[0]
port 11 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 y[1]
port 12 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 y[2]
port 13 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 y[3]
port 14 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 y[4]
port 15 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 y[5]
port 16 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 y[6]
port 17 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 y[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 345014
string GDS_FILE /openlane/designs/lab1/runs/RUN_2025.04.26_11.56.03/results/signoff/lab1.magic.gds
string GDS_START 102522
<< end >>

