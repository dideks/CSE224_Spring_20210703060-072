* NGSPICE file created from lab1.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

.subckt lab1 VGND VPWR x[0] x[1] x[2] x[3] x[4] x[5] x[6] x[7] y[0] y[1] y[2] y[3]
+ y[4] y[5] y[6] y[7]
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput10 net10 VGND VGND VPWR VPWR y[1] sky130_fd_sc_hd__buf_2
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net9 VGND VGND VPWR VPWR y[0] sky130_fd_sc_hd__buf_2
Xoutput11 net11 VGND VGND VPWR VPWR y[2] sky130_fd_sc_hd__buf_2
XFILLER_0_27_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput12 net12 VGND VGND VPWR VPWR y[3] sky130_fd_sc_hd__buf_2
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR y[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_27_ net1 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput14 net14 VGND VGND VPWR VPWR y[5] sky130_fd_sc_hd__buf_2
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_26_ _00_ _09_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__nor2_1
XFILLER_0_21_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR y[6] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_25_ net2 net1 VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput16 net16 VGND VGND VPWR VPWR y[7] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_17_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_24_ net8 _06_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__xor2_1
XFILLER_0_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_47 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23_ _08_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_22_ _06_ _07_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_21_ net5 net6 _02_ net7 VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_20_ net5 net6 net7 _02_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__or4_2
Xinput1 x[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_27_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_11_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 x[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 x[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 x[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_0_14_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 x[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 x[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 x[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 x[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_19_ net6 _04_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18_ _04_ _05_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17_ net5 _02_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16_ net5 _02_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ _03_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14_ _01_ _02_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_9_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13_ net2 net1 net3 net4 VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__or4_4
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12_ net2 net1 net3 net4 VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11_ net3 _00_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10_ net2 net1 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_8_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
.ends

