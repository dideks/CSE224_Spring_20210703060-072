VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lab1
  CLASS BLOCK ;
  FOREIGN lab1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 19.115 10.640 20.715 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.310 10.640 42.910 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 63.505 10.640 65.105 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.700 10.640 87.300 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 22.900 94.540 24.500 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.940 94.540 43.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 60.980 94.540 62.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 80.020 94.540 81.620 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.600 94.540 21.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 38.640 94.540 40.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 57.680 94.540 59.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.720 94.540 78.320 ;
    END
  END VPWR
  PIN x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END x[7]
  PIN y[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END y[0]
  PIN y[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END y[1]
  PIN y[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END y[2]
  PIN y[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END y[3]
  PIN y[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END y[4]
  PIN y[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END y[5]
  PIN y[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END y[6]
  PIN y[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END y[7]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 4.210 10.640 94.300 87.280 ;
      LAYER met2 ;
        RECT 4.230 10.695 92.820 87.225 ;
      LAYER met3 ;
        RECT 3.990 75.840 87.290 87.205 ;
        RECT 4.400 74.440 87.290 75.840 ;
        RECT 3.990 72.440 87.290 74.440 ;
        RECT 4.400 71.040 87.290 72.440 ;
        RECT 3.990 69.040 87.290 71.040 ;
        RECT 4.400 67.640 87.290 69.040 ;
        RECT 3.990 65.640 87.290 67.640 ;
        RECT 4.400 64.240 87.290 65.640 ;
        RECT 3.990 62.240 87.290 64.240 ;
        RECT 4.400 60.840 87.290 62.240 ;
        RECT 3.990 58.840 87.290 60.840 ;
        RECT 4.400 57.440 87.290 58.840 ;
        RECT 3.990 55.440 87.290 57.440 ;
        RECT 4.400 54.040 87.290 55.440 ;
        RECT 3.990 52.040 87.290 54.040 ;
        RECT 4.400 50.640 87.290 52.040 ;
        RECT 3.990 48.640 87.290 50.640 ;
        RECT 4.400 47.240 87.290 48.640 ;
        RECT 3.990 45.240 87.290 47.240 ;
        RECT 4.400 43.840 87.290 45.240 ;
        RECT 3.990 41.840 87.290 43.840 ;
        RECT 4.400 40.440 87.290 41.840 ;
        RECT 3.990 38.440 87.290 40.440 ;
        RECT 4.400 37.040 87.290 38.440 ;
        RECT 3.990 35.040 87.290 37.040 ;
        RECT 4.400 33.640 87.290 35.040 ;
        RECT 3.990 31.640 87.290 33.640 ;
        RECT 4.400 30.240 87.290 31.640 ;
        RECT 3.990 28.240 87.290 30.240 ;
        RECT 4.400 26.840 87.290 28.240 ;
        RECT 3.990 24.840 87.290 26.840 ;
        RECT 4.400 23.440 87.290 24.840 ;
        RECT 3.990 10.715 87.290 23.440 ;
  END
END lab1
END LIBRARY

