magic
tech sky130A
magscale 1 2
timestamp 1745668593
<< checkpaint >>
rect -3932 -1804 22840 21388
<< viali >>
rect 6837 17289 6871 17323
rect 6377 17153 6411 17187
rect 6837 17153 6871 17187
rect 6653 17017 6687 17051
rect 6515 16949 6549 16983
rect 15209 16745 15243 16779
rect 15117 16609 15151 16643
rect 4169 16541 4203 16575
rect 15025 16541 15059 16575
rect 15301 16473 15335 16507
rect 3985 16405 4019 16439
rect 14841 16405 14875 16439
rect 17509 16065 17543 16099
rect 16865 15997 16899 16031
rect 17417 15997 17451 16031
rect 1685 15453 1719 15487
rect 15577 15453 15611 15487
rect 15669 15453 15703 15487
rect 1501 15317 1535 15351
rect 15393 15317 15427 15351
rect 1501 14501 1535 14535
rect 18153 14433 18187 14467
rect 1685 14365 1719 14399
rect 17969 14365 18003 14399
rect 18061 14365 18095 14399
rect 18245 14365 18279 14399
rect 18429 14229 18463 14263
rect 8861 14025 8895 14059
rect 1685 13889 1719 13923
rect 9045 13889 9079 13923
rect 18245 13889 18279 13923
rect 18429 13889 18463 13923
rect 18337 13821 18371 13855
rect 1501 13685 1535 13719
rect 5825 13413 5859 13447
rect 5917 13345 5951 13379
rect 1685 13277 1719 13311
rect 5696 13277 5730 13311
rect 5549 13209 5583 13243
rect 1501 13141 1535 13175
rect 6193 13141 6227 13175
rect 1685 12869 1719 12903
rect 1501 12801 1535 12835
rect 1685 11713 1719 11747
rect 1501 11577 1535 11611
rect 1593 11305 1627 11339
rect 1501 11033 1535 11067
rect 1501 10625 1535 10659
rect 1685 10489 1719 10523
rect 1593 10217 1627 10251
rect 1409 10013 1443 10047
rect 8217 9605 8251 9639
rect 8033 9537 8067 9571
rect 7849 9469 7883 9503
rect 1593 9129 1627 9163
rect 1409 8925 1443 8959
rect 1593 8585 1627 8619
rect 1409 8449 1443 8483
rect 3801 8449 3835 8483
rect 3893 8381 3927 8415
rect 3433 8245 3467 8279
rect 9137 7973 9171 8007
rect 8953 7905 8987 7939
rect 1685 7837 1719 7871
rect 8401 7837 8435 7871
rect 9413 7769 9447 7803
rect 1501 7701 1535 7735
rect 8217 7701 8251 7735
rect 7573 7497 7607 7531
rect 1685 7429 1719 7463
rect 1501 7361 1535 7395
rect 7941 7361 7975 7395
rect 13921 7361 13955 7395
rect 14105 7361 14139 7395
rect 8033 7293 8067 7327
rect 13921 7225 13955 7259
rect 1501 6409 1535 6443
rect 1685 6273 1719 6307
rect 1685 5661 1719 5695
rect 16497 5661 16531 5695
rect 16681 5661 16715 5695
rect 16589 5593 16623 5627
rect 1501 5525 1535 5559
rect 1501 5185 1535 5219
rect 1593 4981 1627 5015
rect 3893 4641 3927 4675
rect 4077 4573 4111 4607
rect 4261 4437 4295 4471
rect 5825 2601 5859 2635
rect 5825 2397 5859 2431
rect 6009 2397 6043 2431
<< metal1 >>
rect 1104 17434 18860 17456
rect 1104 17382 3829 17434
rect 3881 17382 3893 17434
rect 3945 17382 3957 17434
rect 4009 17382 4021 17434
rect 4073 17382 4085 17434
rect 4137 17382 8268 17434
rect 8320 17382 8332 17434
rect 8384 17382 8396 17434
rect 8448 17382 8460 17434
rect 8512 17382 8524 17434
rect 8576 17382 12707 17434
rect 12759 17382 12771 17434
rect 12823 17382 12835 17434
rect 12887 17382 12899 17434
rect 12951 17382 12963 17434
rect 13015 17382 17146 17434
rect 17198 17382 17210 17434
rect 17262 17382 17274 17434
rect 17326 17382 17338 17434
rect 17390 17382 17402 17434
rect 17454 17382 18860 17434
rect 1104 17360 18860 17382
rect 6825 17323 6883 17329
rect 6825 17289 6837 17323
rect 6871 17320 6883 17323
rect 8018 17320 8024 17332
rect 6871 17292 8024 17320
rect 6871 17289 6883 17292
rect 6825 17283 6883 17289
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 15010 17252 15016 17264
rect 6380 17224 15016 17252
rect 6380 17193 6408 17224
rect 15010 17212 15016 17224
rect 15068 17212 15074 17264
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6822 17184 6828 17196
rect 6783 17156 6828 17184
rect 6365 17147 6423 17153
rect 6822 17144 6828 17156
rect 6880 17184 6886 17196
rect 15102 17184 15108 17196
rect 6880 17156 15108 17184
rect 6880 17144 6886 17156
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 6178 17008 6184 17060
rect 6236 17048 6242 17060
rect 6641 17051 6699 17057
rect 6641 17048 6653 17051
rect 6236 17020 6653 17048
rect 6236 17008 6242 17020
rect 6641 17017 6653 17020
rect 6687 17017 6699 17051
rect 6641 17011 6699 17017
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 6503 16983 6561 16989
rect 6503 16980 6515 16983
rect 5408 16952 6515 16980
rect 5408 16940 5414 16952
rect 6503 16949 6515 16952
rect 6549 16980 6561 16983
rect 15194 16980 15200 16992
rect 6549 16952 15200 16980
rect 6549 16949 6561 16952
rect 6503 16943 6561 16949
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 15194 16736 15200 16788
rect 15252 16736 15258 16788
rect 15102 16600 15108 16652
rect 15160 16600 15166 16652
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 5810 16572 5816 16584
rect 4203 16544 5816 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 15010 16532 15016 16584
rect 15068 16532 15074 16584
rect 15286 16464 15292 16516
rect 15344 16464 15350 16516
rect 3602 16396 3608 16448
rect 3660 16436 3666 16448
rect 3973 16439 4031 16445
rect 3973 16436 3985 16439
rect 3660 16408 3985 16436
rect 3660 16396 3666 16408
rect 3973 16405 3985 16408
rect 4019 16405 4031 16439
rect 3973 16399 4031 16405
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 14829 16439 14887 16445
rect 14829 16436 14841 16439
rect 11112 16408 14841 16436
rect 11112 16396 11118 16408
rect 14829 16405 14841 16408
rect 14875 16405 14887 16439
rect 14829 16399 14887 16405
rect 1104 16346 18860 16368
rect 1104 16294 3829 16346
rect 3881 16294 3893 16346
rect 3945 16294 3957 16346
rect 4009 16294 4021 16346
rect 4073 16294 4085 16346
rect 4137 16294 8268 16346
rect 8320 16294 8332 16346
rect 8384 16294 8396 16346
rect 8448 16294 8460 16346
rect 8512 16294 8524 16346
rect 8576 16294 12707 16346
rect 12759 16294 12771 16346
rect 12823 16294 12835 16346
rect 12887 16294 12899 16346
rect 12951 16294 12963 16346
rect 13015 16294 17146 16346
rect 17198 16294 17210 16346
rect 17262 16294 17274 16346
rect 17326 16294 17338 16346
rect 17390 16294 17402 16346
rect 17454 16294 18860 16346
rect 1104 16272 18860 16294
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 17497 16099 17555 16105
rect 17497 16096 17509 16099
rect 15252 16068 17509 16096
rect 15252 16056 15258 16068
rect 17497 16065 17509 16068
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 1820 16000 16865 16028
rect 1820 15988 1826 16000
rect 16853 15997 16865 16000
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 17034 15988 17040 16040
rect 17092 16028 17098 16040
rect 17405 16031 17463 16037
rect 17405 16028 17417 16031
rect 17092 16000 17417 16028
rect 17092 15988 17098 16000
rect 17405 15997 17417 16000
rect 17451 15997 17463 16031
rect 17405 15991 17463 15997
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 1670 15444 1676 15496
rect 1728 15444 1734 15496
rect 6178 15444 6184 15496
rect 6236 15484 6242 15496
rect 15286 15484 15292 15496
rect 6236 15456 15292 15484
rect 6236 15444 6242 15456
rect 15286 15444 15292 15456
rect 15344 15484 15350 15496
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 15344 15456 15577 15484
rect 15344 15444 15350 15456
rect 15565 15453 15577 15456
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 15657 15487 15715 15493
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 14090 15376 14096 15428
rect 14148 15416 14154 15428
rect 15010 15416 15016 15428
rect 14148 15388 15016 15416
rect 14148 15376 14154 15388
rect 15010 15376 15016 15388
rect 15068 15416 15074 15428
rect 15672 15416 15700 15447
rect 15068 15388 15700 15416
rect 15068 15376 15074 15388
rect 1486 15308 1492 15360
rect 1544 15308 1550 15360
rect 15378 15308 15384 15360
rect 15436 15308 15442 15360
rect 1104 15258 18860 15280
rect 1104 15206 3829 15258
rect 3881 15206 3893 15258
rect 3945 15206 3957 15258
rect 4009 15206 4021 15258
rect 4073 15206 4085 15258
rect 4137 15206 8268 15258
rect 8320 15206 8332 15258
rect 8384 15206 8396 15258
rect 8448 15206 8460 15258
rect 8512 15206 8524 15258
rect 8576 15206 12707 15258
rect 12759 15206 12771 15258
rect 12823 15206 12835 15258
rect 12887 15206 12899 15258
rect 12951 15206 12963 15258
rect 13015 15206 17146 15258
rect 17198 15206 17210 15258
rect 17262 15206 17274 15258
rect 17326 15206 17338 15258
rect 17390 15206 17402 15258
rect 17454 15206 18860 15258
rect 1104 15184 18860 15206
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 842 14492 848 14544
rect 900 14532 906 14544
rect 1489 14535 1547 14541
rect 1489 14532 1501 14535
rect 900 14504 1501 14532
rect 900 14492 906 14504
rect 1489 14501 1501 14504
rect 1535 14501 1547 14535
rect 1489 14495 1547 14501
rect 5810 14424 5816 14476
rect 5868 14464 5874 14476
rect 18138 14464 18144 14476
rect 5868 14436 18144 14464
rect 5868 14424 5874 14436
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1854 14396 1860 14408
rect 1719 14368 1860 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17957 14399 18015 14405
rect 17957 14396 17969 14399
rect 17000 14368 17969 14396
rect 17000 14356 17006 14368
rect 17957 14365 17969 14368
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18506 14396 18512 14408
rect 18279 14368 18512 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 18064 14328 18092 14359
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 8168 14300 18092 14328
rect 8168 14288 8174 14300
rect 18414 14220 18420 14272
rect 18472 14220 18478 14272
rect 1104 14170 18860 14192
rect 1104 14118 3829 14170
rect 3881 14118 3893 14170
rect 3945 14118 3957 14170
rect 4009 14118 4021 14170
rect 4073 14118 4085 14170
rect 4137 14118 8268 14170
rect 8320 14118 8332 14170
rect 8384 14118 8396 14170
rect 8448 14118 8460 14170
rect 8512 14118 8524 14170
rect 8576 14118 12707 14170
rect 12759 14118 12771 14170
rect 12823 14118 12835 14170
rect 12887 14118 12899 14170
rect 12951 14118 12963 14170
rect 13015 14118 17146 14170
rect 17198 14118 17210 14170
rect 17262 14118 17274 14170
rect 17326 14118 17338 14170
rect 17390 14118 17402 14170
rect 17454 14118 18860 14170
rect 1104 14096 18860 14118
rect 8849 14059 8907 14065
rect 8849 14056 8861 14059
rect 6886 14028 8861 14056
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 6886 13920 6914 14028
rect 8849 14025 8861 14028
rect 8895 14025 8907 14059
rect 8849 14019 8907 14025
rect 1719 13892 6914 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 9030 13880 9036 13932
rect 9088 13880 9094 13932
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 18196 13892 18245 13920
rect 18196 13880 18202 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13920 18475 13923
rect 18506 13920 18512 13932
rect 18463 13892 18512 13920
rect 18463 13889 18475 13892
rect 18417 13883 18475 13889
rect 18506 13880 18512 13892
rect 18564 13880 18570 13932
rect 17494 13812 17500 13864
rect 17552 13852 17558 13864
rect 18325 13855 18383 13861
rect 18325 13852 18337 13855
rect 17552 13824 18337 13852
rect 17552 13812 17558 13824
rect 18325 13821 18337 13824
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 1486 13676 1492 13728
rect 1544 13676 1550 13728
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 5810 13404 5816 13456
rect 5868 13404 5874 13456
rect 3694 13336 3700 13388
rect 3752 13376 3758 13388
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 3752 13348 5917 13376
rect 3752 13336 3758 13348
rect 5905 13345 5917 13348
rect 5951 13376 5963 13379
rect 18506 13376 18512 13388
rect 5951 13348 18512 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 18506 13336 18512 13348
rect 18564 13336 18570 13388
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 3602 13308 3608 13320
rect 1719 13280 3608 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 3602 13268 3608 13280
rect 3660 13268 3666 13320
rect 5718 13317 5724 13320
rect 5684 13311 5724 13317
rect 5684 13277 5696 13311
rect 5684 13271 5724 13277
rect 5718 13268 5724 13271
rect 5776 13268 5782 13320
rect 4798 13200 4804 13252
rect 4856 13240 4862 13252
rect 5537 13243 5595 13249
rect 5537 13240 5549 13243
rect 4856 13212 5549 13240
rect 4856 13200 4862 13212
rect 5537 13209 5549 13212
rect 5583 13240 5595 13243
rect 16942 13240 16948 13252
rect 5583 13212 16948 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 16942 13200 16948 13212
rect 17000 13200 17006 13252
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1489 13175 1547 13181
rect 1489 13172 1501 13175
rect 900 13144 1501 13172
rect 900 13132 906 13144
rect 1489 13141 1501 13144
rect 1535 13141 1547 13175
rect 1489 13135 1547 13141
rect 6178 13132 6184 13184
rect 6236 13132 6242 13184
rect 1104 13082 18860 13104
rect 1104 13030 3829 13082
rect 3881 13030 3893 13082
rect 3945 13030 3957 13082
rect 4009 13030 4021 13082
rect 4073 13030 4085 13082
rect 4137 13030 8268 13082
rect 8320 13030 8332 13082
rect 8384 13030 8396 13082
rect 8448 13030 8460 13082
rect 8512 13030 8524 13082
rect 8576 13030 12707 13082
rect 12759 13030 12771 13082
rect 12823 13030 12835 13082
rect 12887 13030 12899 13082
rect 12951 13030 12963 13082
rect 13015 13030 17146 13082
rect 17198 13030 17210 13082
rect 17262 13030 17274 13082
rect 17326 13030 17338 13082
rect 17390 13030 17402 13082
rect 17454 13030 18860 13082
rect 1104 13008 18860 13030
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 5350 12900 5356 12912
rect 1719 12872 5356 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 1486 12792 1492 12844
rect 1544 12792 1550 12844
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 1104 11994 18860 12016
rect 1104 11942 3829 11994
rect 3881 11942 3893 11994
rect 3945 11942 3957 11994
rect 4009 11942 4021 11994
rect 4073 11942 4085 11994
rect 4137 11942 8268 11994
rect 8320 11942 8332 11994
rect 8384 11942 8396 11994
rect 8448 11942 8460 11994
rect 8512 11942 8524 11994
rect 8576 11942 12707 11994
rect 12759 11942 12771 11994
rect 12823 11942 12835 11994
rect 12887 11942 12899 11994
rect 12951 11942 12963 11994
rect 13015 11942 17146 11994
rect 17198 11942 17210 11994
rect 17262 11942 17274 11994
rect 17326 11942 17338 11994
rect 17390 11942 17402 11994
rect 17454 11942 18860 11994
rect 1104 11920 18860 11942
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 3694 11744 3700 11756
rect 1719 11716 3700 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 842 11568 848 11620
rect 900 11608 906 11620
rect 1489 11611 1547 11617
rect 1489 11608 1501 11611
rect 900 11580 1501 11608
rect 900 11568 906 11580
rect 1489 11577 1501 11580
rect 1535 11577 1547 11611
rect 1489 11571 1547 11577
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 5718 11336 5724 11348
rect 1627 11308 5724 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 5718 11296 5724 11308
rect 5776 11336 5782 11348
rect 8110 11336 8116 11348
rect 5776 11308 8116 11336
rect 5776 11296 5782 11308
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 1486 11024 1492 11076
rect 1544 11024 1550 11076
rect 1104 10906 18860 10928
rect 1104 10854 3829 10906
rect 3881 10854 3893 10906
rect 3945 10854 3957 10906
rect 4009 10854 4021 10906
rect 4073 10854 4085 10906
rect 4137 10854 8268 10906
rect 8320 10854 8332 10906
rect 8384 10854 8396 10906
rect 8448 10854 8460 10906
rect 8512 10854 8524 10906
rect 8576 10854 12707 10906
rect 12759 10854 12771 10906
rect 12823 10854 12835 10906
rect 12887 10854 12899 10906
rect 12951 10854 12963 10906
rect 13015 10854 17146 10906
rect 17198 10854 17210 10906
rect 17262 10854 17274 10906
rect 17326 10854 17338 10906
rect 17390 10854 17402 10906
rect 17454 10854 18860 10906
rect 1104 10832 18860 10854
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 1489 10659 1547 10665
rect 1489 10656 1501 10659
rect 900 10628 1501 10656
rect 900 10616 906 10628
rect 1489 10625 1501 10628
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10520 1731 10523
rect 3602 10520 3608 10532
rect 1719 10492 3608 10520
rect 1719 10489 1731 10492
rect 1673 10483 1731 10489
rect 3602 10480 3608 10492
rect 3660 10480 3666 10532
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 4798 10248 4804 10260
rect 1627 10220 4804 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1104 9818 18860 9840
rect 1104 9766 3829 9818
rect 3881 9766 3893 9818
rect 3945 9766 3957 9818
rect 4009 9766 4021 9818
rect 4073 9766 4085 9818
rect 4137 9766 8268 9818
rect 8320 9766 8332 9818
rect 8384 9766 8396 9818
rect 8448 9766 8460 9818
rect 8512 9766 8524 9818
rect 8576 9766 12707 9818
rect 12759 9766 12771 9818
rect 12823 9766 12835 9818
rect 12887 9766 12899 9818
rect 12951 9766 12963 9818
rect 13015 9766 17146 9818
rect 17198 9766 17210 9818
rect 17262 9766 17274 9818
rect 17326 9766 17338 9818
rect 17390 9766 17402 9818
rect 17454 9766 18860 9818
rect 1104 9744 18860 9766
rect 8205 9639 8263 9645
rect 8205 9605 8217 9639
rect 8251 9636 8263 9639
rect 9030 9636 9036 9648
rect 8251 9608 9036 9636
rect 8251 9605 8263 9608
rect 8205 9599 8263 9605
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 8018 9528 8024 9580
rect 8076 9528 8082 9580
rect 7466 9460 7472 9512
rect 7524 9500 7530 9512
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 7524 9472 7849 9500
rect 7524 9460 7530 9472
rect 7837 9469 7849 9472
rect 7883 9500 7895 9503
rect 11054 9500 11060 9512
rect 7883 9472 11060 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 6822 9160 6828 9172
rect 1627 9132 6828 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1104 8730 18860 8752
rect 1104 8678 3829 8730
rect 3881 8678 3893 8730
rect 3945 8678 3957 8730
rect 4009 8678 4021 8730
rect 4073 8678 4085 8730
rect 4137 8678 8268 8730
rect 8320 8678 8332 8730
rect 8384 8678 8396 8730
rect 8448 8678 8460 8730
rect 8512 8678 8524 8730
rect 8576 8678 12707 8730
rect 12759 8678 12771 8730
rect 12823 8678 12835 8730
rect 12887 8678 12899 8730
rect 12951 8678 12963 8730
rect 13015 8678 17146 8730
rect 17198 8678 17210 8730
rect 17262 8678 17274 8730
rect 17326 8678 17338 8730
rect 17390 8678 17402 8730
rect 17454 8678 18860 8730
rect 1104 8656 18860 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1596 8480 1624 8579
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 1596 8452 3801 8480
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 3881 8415 3939 8421
rect 3881 8381 3893 8415
rect 3927 8412 3939 8415
rect 7466 8412 7472 8424
rect 3927 8384 7472 8412
rect 3927 8381 3939 8384
rect 3881 8375 3939 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 2832 8248 3433 8276
rect 2832 8236 2838 8248
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 6178 7964 6184 8016
rect 6236 8004 6242 8016
rect 9122 8004 9128 8016
rect 6236 7976 9128 8004
rect 6236 7964 6242 7976
rect 9122 7964 9128 7976
rect 9180 7964 9186 8016
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8404 7908 8953 7936
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2774 7868 2780 7880
rect 1719 7840 2780 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 8404 7877 8432 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 9401 7803 9459 7809
rect 9401 7769 9413 7803
rect 9447 7800 9459 7803
rect 18414 7800 18420 7812
rect 9447 7772 18420 7800
rect 9447 7769 9459 7772
rect 9401 7763 9459 7769
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 842 7692 848 7744
rect 900 7732 906 7744
rect 1489 7735 1547 7741
rect 1489 7732 1501 7735
rect 900 7704 1501 7732
rect 900 7692 906 7704
rect 1489 7701 1501 7704
rect 1535 7701 1547 7735
rect 1489 7695 1547 7701
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 6972 7704 8217 7732
rect 6972 7692 6978 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 1104 7642 18860 7664
rect 1104 7590 3829 7642
rect 3881 7590 3893 7642
rect 3945 7590 3957 7642
rect 4009 7590 4021 7642
rect 4073 7590 4085 7642
rect 4137 7590 8268 7642
rect 8320 7590 8332 7642
rect 8384 7590 8396 7642
rect 8448 7590 8460 7642
rect 8512 7590 8524 7642
rect 8576 7590 12707 7642
rect 12759 7590 12771 7642
rect 12823 7590 12835 7642
rect 12887 7590 12899 7642
rect 12951 7590 12963 7642
rect 13015 7590 17146 7642
rect 17198 7590 17210 7642
rect 17262 7590 17274 7642
rect 17326 7590 17338 7642
rect 17390 7590 17402 7642
rect 17454 7590 18860 7642
rect 1104 7568 18860 7590
rect 3694 7488 3700 7540
rect 3752 7528 3758 7540
rect 7561 7531 7619 7537
rect 7561 7528 7573 7531
rect 3752 7500 7573 7528
rect 3752 7488 3758 7500
rect 7561 7497 7573 7500
rect 7607 7497 7619 7531
rect 7561 7491 7619 7497
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 1719 7432 14044 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8110 7392 8116 7404
rect 7975 7364 8116 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 9122 7352 9128 7404
rect 9180 7392 9186 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 9180 7364 13921 7392
rect 9180 7352 9186 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 14016 7392 14044 7432
rect 14090 7392 14096 7404
rect 14016 7364 14096 7392
rect 13909 7355 13967 7361
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 17494 7324 17500 7336
rect 8067 7296 17500 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 17494 7284 17500 7296
rect 17552 7284 17558 7336
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 17034 7256 17040 7268
rect 13964 7228 17040 7256
rect 13964 7216 13970 7228
rect 17034 7216 17040 7228
rect 17092 7216 17098 7268
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 1104 6554 18860 6576
rect 1104 6502 3829 6554
rect 3881 6502 3893 6554
rect 3945 6502 3957 6554
rect 4009 6502 4021 6554
rect 4073 6502 4085 6554
rect 4137 6502 8268 6554
rect 8320 6502 8332 6554
rect 8384 6502 8396 6554
rect 8448 6502 8460 6554
rect 8512 6502 8524 6554
rect 8576 6502 12707 6554
rect 12759 6502 12771 6554
rect 12823 6502 12835 6554
rect 12887 6502 12899 6554
rect 12951 6502 12963 6554
rect 13015 6502 17146 6554
rect 17198 6502 17210 6554
rect 17262 6502 17274 6554
rect 17326 6502 17338 6554
rect 17390 6502 17402 6554
rect 17454 6502 18860 6554
rect 1104 6480 18860 6502
rect 842 6400 848 6452
rect 900 6440 906 6452
rect 1489 6443 1547 6449
rect 1489 6440 1501 6443
rect 900 6412 1501 6440
rect 900 6400 906 6412
rect 1489 6409 1501 6412
rect 1535 6409 1547 6443
rect 1489 6403 1547 6409
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 1762 6304 1768 6316
rect 1719 6276 1768 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 6914 5692 6920 5704
rect 1719 5664 6920 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 16485 5695 16543 5701
rect 16485 5692 16497 5695
rect 13872 5664 16497 5692
rect 13872 5652 13878 5664
rect 16485 5661 16497 5664
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5692 16727 5695
rect 17494 5692 17500 5704
rect 16715 5664 17500 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 1854 5584 1860 5636
rect 1912 5624 1918 5636
rect 16577 5627 16635 5633
rect 16577 5624 16589 5627
rect 1912 5596 16589 5624
rect 1912 5584 1918 5596
rect 16577 5593 16589 5596
rect 16623 5593 16635 5627
rect 16577 5587 16635 5593
rect 1486 5516 1492 5568
rect 1544 5516 1550 5568
rect 1104 5466 18860 5488
rect 1104 5414 3829 5466
rect 3881 5414 3893 5466
rect 3945 5414 3957 5466
rect 4009 5414 4021 5466
rect 4073 5414 4085 5466
rect 4137 5414 8268 5466
rect 8320 5414 8332 5466
rect 8384 5414 8396 5466
rect 8448 5414 8460 5466
rect 8512 5414 8524 5466
rect 8576 5414 12707 5466
rect 12759 5414 12771 5466
rect 12823 5414 12835 5466
rect 12887 5414 12899 5466
rect 12951 5414 12963 5466
rect 13015 5414 17146 5466
rect 17198 5414 17210 5466
rect 17262 5414 17274 5466
rect 17326 5414 17338 5466
rect 17390 5414 17402 5466
rect 17454 5414 18860 5466
rect 1104 5392 18860 5414
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 900 5188 1501 5216
rect 900 5176 906 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 3694 4632 3700 4684
rect 3752 4672 3758 4684
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 3752 4644 3893 4672
rect 3752 4632 3758 4644
rect 3881 4641 3893 4644
rect 3927 4641 3939 4675
rect 3881 4635 3939 4641
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 1636 4576 4077 4604
rect 1636 4564 1642 4576
rect 4065 4573 4077 4576
rect 4111 4604 4123 4607
rect 5810 4604 5816 4616
rect 4111 4576 5816 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 13814 4468 13820 4480
rect 4295 4440 13820 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 1104 4378 18860 4400
rect 1104 4326 3829 4378
rect 3881 4326 3893 4378
rect 3945 4326 3957 4378
rect 4009 4326 4021 4378
rect 4073 4326 4085 4378
rect 4137 4326 8268 4378
rect 8320 4326 8332 4378
rect 8384 4326 8396 4378
rect 8448 4326 8460 4378
rect 8512 4326 8524 4378
rect 8576 4326 12707 4378
rect 12759 4326 12771 4378
rect 12823 4326 12835 4378
rect 12887 4326 12899 4378
rect 12951 4326 12963 4378
rect 13015 4326 17146 4378
rect 17198 4326 17210 4378
rect 17262 4326 17274 4378
rect 17326 4326 17338 4378
rect 17390 4326 17402 4378
rect 17454 4326 18860 4378
rect 1104 4304 18860 4326
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 1104 3290 18860 3312
rect 1104 3238 3829 3290
rect 3881 3238 3893 3290
rect 3945 3238 3957 3290
rect 4009 3238 4021 3290
rect 4073 3238 4085 3290
rect 4137 3238 8268 3290
rect 8320 3238 8332 3290
rect 8384 3238 8396 3290
rect 8448 3238 8460 3290
rect 8512 3238 8524 3290
rect 8576 3238 12707 3290
rect 12759 3238 12771 3290
rect 12823 3238 12835 3290
rect 12887 3238 12899 3290
rect 12951 3238 12963 3290
rect 13015 3238 17146 3290
rect 17198 3238 17210 3290
rect 17262 3238 17274 3290
rect 17326 3238 17338 3290
rect 17390 3238 17402 3290
rect 17454 3238 18860 3290
rect 1104 3216 18860 3238
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 1728 2604 5825 2632
rect 1728 2592 1734 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 5813 2595 5871 2601
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 13906 2428 13912 2440
rect 6043 2400 13912 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 5828 2360 5856 2391
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 15378 2360 15384 2372
rect 5828 2332 15384 2360
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 1104 2202 18860 2224
rect 1104 2150 3829 2202
rect 3881 2150 3893 2202
rect 3945 2150 3957 2202
rect 4009 2150 4021 2202
rect 4073 2150 4085 2202
rect 4137 2150 8268 2202
rect 8320 2150 8332 2202
rect 8384 2150 8396 2202
rect 8448 2150 8460 2202
rect 8512 2150 8524 2202
rect 8576 2150 12707 2202
rect 12759 2150 12771 2202
rect 12823 2150 12835 2202
rect 12887 2150 12899 2202
rect 12951 2150 12963 2202
rect 13015 2150 17146 2202
rect 17198 2150 17210 2202
rect 17262 2150 17274 2202
rect 17326 2150 17338 2202
rect 17390 2150 17402 2202
rect 17454 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 3829 17382 3881 17434
rect 3893 17382 3945 17434
rect 3957 17382 4009 17434
rect 4021 17382 4073 17434
rect 4085 17382 4137 17434
rect 8268 17382 8320 17434
rect 8332 17382 8384 17434
rect 8396 17382 8448 17434
rect 8460 17382 8512 17434
rect 8524 17382 8576 17434
rect 12707 17382 12759 17434
rect 12771 17382 12823 17434
rect 12835 17382 12887 17434
rect 12899 17382 12951 17434
rect 12963 17382 13015 17434
rect 17146 17382 17198 17434
rect 17210 17382 17262 17434
rect 17274 17382 17326 17434
rect 17338 17382 17390 17434
rect 17402 17382 17454 17434
rect 8024 17280 8076 17332
rect 15016 17212 15068 17264
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 15108 17144 15160 17196
rect 6184 17008 6236 17060
rect 5356 16940 5408 16992
rect 15200 16940 15252 16992
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 15200 16779 15252 16788
rect 15200 16745 15209 16779
rect 15209 16745 15243 16779
rect 15243 16745 15252 16779
rect 15200 16736 15252 16745
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 5816 16532 5868 16584
rect 15016 16575 15068 16584
rect 15016 16541 15025 16575
rect 15025 16541 15059 16575
rect 15059 16541 15068 16575
rect 15016 16532 15068 16541
rect 15292 16507 15344 16516
rect 15292 16473 15301 16507
rect 15301 16473 15335 16507
rect 15335 16473 15344 16507
rect 15292 16464 15344 16473
rect 3608 16396 3660 16448
rect 11060 16396 11112 16448
rect 3829 16294 3881 16346
rect 3893 16294 3945 16346
rect 3957 16294 4009 16346
rect 4021 16294 4073 16346
rect 4085 16294 4137 16346
rect 8268 16294 8320 16346
rect 8332 16294 8384 16346
rect 8396 16294 8448 16346
rect 8460 16294 8512 16346
rect 8524 16294 8576 16346
rect 12707 16294 12759 16346
rect 12771 16294 12823 16346
rect 12835 16294 12887 16346
rect 12899 16294 12951 16346
rect 12963 16294 13015 16346
rect 17146 16294 17198 16346
rect 17210 16294 17262 16346
rect 17274 16294 17326 16346
rect 17338 16294 17390 16346
rect 17402 16294 17454 16346
rect 15200 16056 15252 16108
rect 1768 15988 1820 16040
rect 17040 15988 17092 16040
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 6184 15444 6236 15496
rect 15292 15444 15344 15496
rect 14096 15376 14148 15428
rect 15016 15376 15068 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 3829 15206 3881 15258
rect 3893 15206 3945 15258
rect 3957 15206 4009 15258
rect 4021 15206 4073 15258
rect 4085 15206 4137 15258
rect 8268 15206 8320 15258
rect 8332 15206 8384 15258
rect 8396 15206 8448 15258
rect 8460 15206 8512 15258
rect 8524 15206 8576 15258
rect 12707 15206 12759 15258
rect 12771 15206 12823 15258
rect 12835 15206 12887 15258
rect 12899 15206 12951 15258
rect 12963 15206 13015 15258
rect 17146 15206 17198 15258
rect 17210 15206 17262 15258
rect 17274 15206 17326 15258
rect 17338 15206 17390 15258
rect 17402 15206 17454 15258
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 848 14492 900 14544
rect 5816 14424 5868 14476
rect 18144 14467 18196 14476
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 1860 14356 1912 14408
rect 16948 14356 17000 14408
rect 8116 14288 8168 14340
rect 18512 14356 18564 14408
rect 18420 14263 18472 14272
rect 18420 14229 18429 14263
rect 18429 14229 18463 14263
rect 18463 14229 18472 14263
rect 18420 14220 18472 14229
rect 3829 14118 3881 14170
rect 3893 14118 3945 14170
rect 3957 14118 4009 14170
rect 4021 14118 4073 14170
rect 4085 14118 4137 14170
rect 8268 14118 8320 14170
rect 8332 14118 8384 14170
rect 8396 14118 8448 14170
rect 8460 14118 8512 14170
rect 8524 14118 8576 14170
rect 12707 14118 12759 14170
rect 12771 14118 12823 14170
rect 12835 14118 12887 14170
rect 12899 14118 12951 14170
rect 12963 14118 13015 14170
rect 17146 14118 17198 14170
rect 17210 14118 17262 14170
rect 17274 14118 17326 14170
rect 17338 14118 17390 14170
rect 17402 14118 17454 14170
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 18144 13880 18196 13932
rect 18512 13880 18564 13932
rect 17500 13812 17552 13864
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 5816 13447 5868 13456
rect 5816 13413 5825 13447
rect 5825 13413 5859 13447
rect 5859 13413 5868 13447
rect 5816 13404 5868 13413
rect 3700 13336 3752 13388
rect 18512 13336 18564 13388
rect 3608 13268 3660 13320
rect 5724 13311 5776 13320
rect 5724 13277 5730 13311
rect 5730 13277 5776 13311
rect 5724 13268 5776 13277
rect 4804 13200 4856 13252
rect 16948 13200 17000 13252
rect 848 13132 900 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 3829 13030 3881 13082
rect 3893 13030 3945 13082
rect 3957 13030 4009 13082
rect 4021 13030 4073 13082
rect 4085 13030 4137 13082
rect 8268 13030 8320 13082
rect 8332 13030 8384 13082
rect 8396 13030 8448 13082
rect 8460 13030 8512 13082
rect 8524 13030 8576 13082
rect 12707 13030 12759 13082
rect 12771 13030 12823 13082
rect 12835 13030 12887 13082
rect 12899 13030 12951 13082
rect 12963 13030 13015 13082
rect 17146 13030 17198 13082
rect 17210 13030 17262 13082
rect 17274 13030 17326 13082
rect 17338 13030 17390 13082
rect 17402 13030 17454 13082
rect 5356 12860 5408 12912
rect 1492 12835 1544 12844
rect 1492 12801 1501 12835
rect 1501 12801 1535 12835
rect 1535 12801 1544 12835
rect 1492 12792 1544 12801
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 3829 11942 3881 11994
rect 3893 11942 3945 11994
rect 3957 11942 4009 11994
rect 4021 11942 4073 11994
rect 4085 11942 4137 11994
rect 8268 11942 8320 11994
rect 8332 11942 8384 11994
rect 8396 11942 8448 11994
rect 8460 11942 8512 11994
rect 8524 11942 8576 11994
rect 12707 11942 12759 11994
rect 12771 11942 12823 11994
rect 12835 11942 12887 11994
rect 12899 11942 12951 11994
rect 12963 11942 13015 11994
rect 17146 11942 17198 11994
rect 17210 11942 17262 11994
rect 17274 11942 17326 11994
rect 17338 11942 17390 11994
rect 17402 11942 17454 11994
rect 3700 11704 3752 11756
rect 848 11568 900 11620
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 5724 11296 5776 11348
rect 8116 11296 8168 11348
rect 1492 11067 1544 11076
rect 1492 11033 1501 11067
rect 1501 11033 1535 11067
rect 1535 11033 1544 11067
rect 1492 11024 1544 11033
rect 3829 10854 3881 10906
rect 3893 10854 3945 10906
rect 3957 10854 4009 10906
rect 4021 10854 4073 10906
rect 4085 10854 4137 10906
rect 8268 10854 8320 10906
rect 8332 10854 8384 10906
rect 8396 10854 8448 10906
rect 8460 10854 8512 10906
rect 8524 10854 8576 10906
rect 12707 10854 12759 10906
rect 12771 10854 12823 10906
rect 12835 10854 12887 10906
rect 12899 10854 12951 10906
rect 12963 10854 13015 10906
rect 17146 10854 17198 10906
rect 17210 10854 17262 10906
rect 17274 10854 17326 10906
rect 17338 10854 17390 10906
rect 17402 10854 17454 10906
rect 848 10616 900 10668
rect 3608 10480 3660 10532
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 4804 10208 4856 10260
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3829 9766 3881 9818
rect 3893 9766 3945 9818
rect 3957 9766 4009 9818
rect 4021 9766 4073 9818
rect 4085 9766 4137 9818
rect 8268 9766 8320 9818
rect 8332 9766 8384 9818
rect 8396 9766 8448 9818
rect 8460 9766 8512 9818
rect 8524 9766 8576 9818
rect 12707 9766 12759 9818
rect 12771 9766 12823 9818
rect 12835 9766 12887 9818
rect 12899 9766 12951 9818
rect 12963 9766 13015 9818
rect 17146 9766 17198 9818
rect 17210 9766 17262 9818
rect 17274 9766 17326 9818
rect 17338 9766 17390 9818
rect 17402 9766 17454 9818
rect 9036 9596 9088 9648
rect 8024 9571 8076 9580
rect 8024 9537 8033 9571
rect 8033 9537 8067 9571
rect 8067 9537 8076 9571
rect 8024 9528 8076 9537
rect 7472 9460 7524 9512
rect 11060 9460 11112 9512
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 6828 9120 6880 9172
rect 848 8916 900 8968
rect 3829 8678 3881 8730
rect 3893 8678 3945 8730
rect 3957 8678 4009 8730
rect 4021 8678 4073 8730
rect 4085 8678 4137 8730
rect 8268 8678 8320 8730
rect 8332 8678 8384 8730
rect 8396 8678 8448 8730
rect 8460 8678 8512 8730
rect 8524 8678 8576 8730
rect 12707 8678 12759 8730
rect 12771 8678 12823 8730
rect 12835 8678 12887 8730
rect 12899 8678 12951 8730
rect 12963 8678 13015 8730
rect 17146 8678 17198 8730
rect 17210 8678 17262 8730
rect 17274 8678 17326 8730
rect 17338 8678 17390 8730
rect 17402 8678 17454 8730
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 7472 8372 7524 8424
rect 2780 8236 2832 8288
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 6184 7964 6236 8016
rect 9128 8007 9180 8016
rect 9128 7973 9137 8007
rect 9137 7973 9171 8007
rect 9171 7973 9180 8007
rect 9128 7964 9180 7973
rect 2780 7828 2832 7880
rect 18420 7760 18472 7812
rect 848 7692 900 7744
rect 6920 7692 6972 7744
rect 3829 7590 3881 7642
rect 3893 7590 3945 7642
rect 3957 7590 4009 7642
rect 4021 7590 4073 7642
rect 4085 7590 4137 7642
rect 8268 7590 8320 7642
rect 8332 7590 8384 7642
rect 8396 7590 8448 7642
rect 8460 7590 8512 7642
rect 8524 7590 8576 7642
rect 12707 7590 12759 7642
rect 12771 7590 12823 7642
rect 12835 7590 12887 7642
rect 12899 7590 12951 7642
rect 12963 7590 13015 7642
rect 17146 7590 17198 7642
rect 17210 7590 17262 7642
rect 17274 7590 17326 7642
rect 17338 7590 17390 7642
rect 17402 7590 17454 7642
rect 3700 7488 3752 7540
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 8116 7352 8168 7404
rect 9128 7352 9180 7404
rect 14096 7395 14148 7404
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 17500 7284 17552 7336
rect 13912 7259 13964 7268
rect 13912 7225 13921 7259
rect 13921 7225 13955 7259
rect 13955 7225 13964 7259
rect 13912 7216 13964 7225
rect 17040 7216 17092 7268
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 3829 6502 3881 6554
rect 3893 6502 3945 6554
rect 3957 6502 4009 6554
rect 4021 6502 4073 6554
rect 4085 6502 4137 6554
rect 8268 6502 8320 6554
rect 8332 6502 8384 6554
rect 8396 6502 8448 6554
rect 8460 6502 8512 6554
rect 8524 6502 8576 6554
rect 12707 6502 12759 6554
rect 12771 6502 12823 6554
rect 12835 6502 12887 6554
rect 12899 6502 12951 6554
rect 12963 6502 13015 6554
rect 17146 6502 17198 6554
rect 17210 6502 17262 6554
rect 17274 6502 17326 6554
rect 17338 6502 17390 6554
rect 17402 6502 17454 6554
rect 848 6400 900 6452
rect 1768 6264 1820 6316
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 6920 5652 6972 5704
rect 13820 5652 13872 5704
rect 17500 5652 17552 5704
rect 1860 5584 1912 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 3829 5414 3881 5466
rect 3893 5414 3945 5466
rect 3957 5414 4009 5466
rect 4021 5414 4073 5466
rect 4085 5414 4137 5466
rect 8268 5414 8320 5466
rect 8332 5414 8384 5466
rect 8396 5414 8448 5466
rect 8460 5414 8512 5466
rect 8524 5414 8576 5466
rect 12707 5414 12759 5466
rect 12771 5414 12823 5466
rect 12835 5414 12887 5466
rect 12899 5414 12951 5466
rect 12963 5414 13015 5466
rect 17146 5414 17198 5466
rect 17210 5414 17262 5466
rect 17274 5414 17326 5466
rect 17338 5414 17390 5466
rect 17402 5414 17454 5466
rect 848 5176 900 5228
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 3700 4632 3752 4684
rect 1584 4564 1636 4616
rect 5816 4564 5868 4616
rect 13820 4428 13872 4480
rect 3829 4326 3881 4378
rect 3893 4326 3945 4378
rect 3957 4326 4009 4378
rect 4021 4326 4073 4378
rect 4085 4326 4137 4378
rect 8268 4326 8320 4378
rect 8332 4326 8384 4378
rect 8396 4326 8448 4378
rect 8460 4326 8512 4378
rect 8524 4326 8576 4378
rect 12707 4326 12759 4378
rect 12771 4326 12823 4378
rect 12835 4326 12887 4378
rect 12899 4326 12951 4378
rect 12963 4326 13015 4378
rect 17146 4326 17198 4378
rect 17210 4326 17262 4378
rect 17274 4326 17326 4378
rect 17338 4326 17390 4378
rect 17402 4326 17454 4378
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 3829 3238 3881 3290
rect 3893 3238 3945 3290
rect 3957 3238 4009 3290
rect 4021 3238 4073 3290
rect 4085 3238 4137 3290
rect 8268 3238 8320 3290
rect 8332 3238 8384 3290
rect 8396 3238 8448 3290
rect 8460 3238 8512 3290
rect 8524 3238 8576 3290
rect 12707 3238 12759 3290
rect 12771 3238 12823 3290
rect 12835 3238 12887 3290
rect 12899 3238 12951 3290
rect 12963 3238 13015 3290
rect 17146 3238 17198 3290
rect 17210 3238 17262 3290
rect 17274 3238 17326 3290
rect 17338 3238 17390 3290
rect 17402 3238 17454 3290
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 1676 2592 1728 2644
rect 13912 2388 13964 2440
rect 15384 2320 15436 2372
rect 3829 2150 3881 2202
rect 3893 2150 3945 2202
rect 3957 2150 4009 2202
rect 4021 2150 4073 2202
rect 4085 2150 4137 2202
rect 8268 2150 8320 2202
rect 8332 2150 8384 2202
rect 8396 2150 8448 2202
rect 8460 2150 8512 2202
rect 8524 2150 8576 2202
rect 12707 2150 12759 2202
rect 12771 2150 12823 2202
rect 12835 2150 12887 2202
rect 12899 2150 12951 2202
rect 12963 2150 13015 2202
rect 17146 2150 17198 2202
rect 17210 2150 17262 2202
rect 17274 2150 17326 2202
rect 17338 2150 17390 2202
rect 17402 2150 17454 2202
<< metal2 >>
rect 3829 17436 4137 17445
rect 3829 17434 3835 17436
rect 3891 17434 3915 17436
rect 3971 17434 3995 17436
rect 4051 17434 4075 17436
rect 4131 17434 4137 17436
rect 3891 17382 3893 17434
rect 4073 17382 4075 17434
rect 3829 17380 3835 17382
rect 3891 17380 3915 17382
rect 3971 17380 3995 17382
rect 4051 17380 4075 17382
rect 4131 17380 4137 17382
rect 3829 17371 4137 17380
rect 8268 17436 8576 17445
rect 8268 17434 8274 17436
rect 8330 17434 8354 17436
rect 8410 17434 8434 17436
rect 8490 17434 8514 17436
rect 8570 17434 8576 17436
rect 8330 17382 8332 17434
rect 8512 17382 8514 17434
rect 8268 17380 8274 17382
rect 8330 17380 8354 17382
rect 8410 17380 8434 17382
rect 8490 17380 8514 17382
rect 8570 17380 8576 17382
rect 8268 17371 8576 17380
rect 12707 17436 13015 17445
rect 12707 17434 12713 17436
rect 12769 17434 12793 17436
rect 12849 17434 12873 17436
rect 12929 17434 12953 17436
rect 13009 17434 13015 17436
rect 12769 17382 12771 17434
rect 12951 17382 12953 17434
rect 12707 17380 12713 17382
rect 12769 17380 12793 17382
rect 12849 17380 12873 17382
rect 12929 17380 12953 17382
rect 13009 17380 13015 17382
rect 12707 17371 13015 17380
rect 17146 17436 17454 17445
rect 17146 17434 17152 17436
rect 17208 17434 17232 17436
rect 17288 17434 17312 17436
rect 17368 17434 17392 17436
rect 17448 17434 17454 17436
rect 17208 17382 17210 17434
rect 17390 17382 17392 17434
rect 17146 17380 17152 17382
rect 17208 17380 17232 17382
rect 17288 17380 17312 17382
rect 17368 17380 17392 17382
rect 17448 17380 17454 17382
rect 17146 17371 17454 17380
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15065 1532 15302
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 848 14544 900 14550
rect 846 14512 848 14521
rect 900 14512 902 14521
rect 846 14447 902 14456
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 1544 13696 1546 13705
rect 1490 13631 1546 13640
rect 848 13184 900 13190
rect 846 13152 848 13161
rect 900 13152 902 13161
rect 846 13087 902 13096
rect 1492 12844 1544 12850
rect 1492 12786 1544 12792
rect 1504 12345 1532 12786
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 848 11620 900 11626
rect 848 11562 900 11568
rect 860 11529 888 11562
rect 846 11520 902 11529
rect 846 11455 902 11464
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1504 10985 1532 11018
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 860 10441 888 10610
rect 846 10432 902 10441
rect 846 10367 902 10376
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 846 9072 902 9081
rect 846 9007 902 9016
rect 860 8974 888 9007
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 848 7744 900 7750
rect 846 7712 848 7721
rect 900 7712 902 7721
rect 846 7647 902 7656
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6905 1532 7346
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 848 6452 900 6458
rect 848 6394 900 6400
rect 860 6361 888 6394
rect 846 6352 902 6361
rect 846 6287 902 6296
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 1584 5024 1636 5030
rect 846 4992 902 5001
rect 1584 4966 1636 4972
rect 846 4927 902 4936
rect 1596 4622 1624 4966
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1688 2650 1716 15438
rect 1780 6322 1808 15982
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1872 5642 1900 14350
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 3620 13326 3648 16390
rect 3829 16348 4137 16357
rect 3829 16346 3835 16348
rect 3891 16346 3915 16348
rect 3971 16346 3995 16348
rect 4051 16346 4075 16348
rect 4131 16346 4137 16348
rect 3891 16294 3893 16346
rect 4073 16294 4075 16346
rect 3829 16292 3835 16294
rect 3891 16292 3915 16294
rect 3971 16292 3995 16294
rect 4051 16292 4075 16294
rect 4131 16292 4137 16294
rect 3829 16283 4137 16292
rect 3829 15260 4137 15269
rect 3829 15258 3835 15260
rect 3891 15258 3915 15260
rect 3971 15258 3995 15260
rect 4051 15258 4075 15260
rect 4131 15258 4137 15260
rect 3891 15206 3893 15258
rect 4073 15206 4075 15258
rect 3829 15204 3835 15206
rect 3891 15204 3915 15206
rect 3971 15204 3995 15206
rect 4051 15204 4075 15206
rect 4131 15204 4137 15206
rect 3829 15195 4137 15204
rect 3829 14172 4137 14181
rect 3829 14170 3835 14172
rect 3891 14170 3915 14172
rect 3971 14170 3995 14172
rect 4051 14170 4075 14172
rect 4131 14170 4137 14172
rect 3891 14118 3893 14170
rect 4073 14118 4075 14170
rect 3829 14116 3835 14118
rect 3891 14116 3915 14118
rect 3971 14116 3995 14118
rect 4051 14116 4075 14118
rect 4131 14116 4137 14118
rect 3829 14107 4137 14116
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3608 13320 3660 13326
rect 3608 13262 3660 13268
rect 3712 13138 3740 13330
rect 4804 13252 4856 13258
rect 4804 13194 4856 13200
rect 3620 13110 3740 13138
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 3620 10538 3648 13110
rect 3829 13084 4137 13093
rect 3829 13082 3835 13084
rect 3891 13082 3915 13084
rect 3971 13082 3995 13084
rect 4051 13082 4075 13084
rect 4131 13082 4137 13084
rect 3891 13030 3893 13082
rect 4073 13030 4075 13082
rect 3829 13028 3835 13030
rect 3891 13028 3915 13030
rect 3971 13028 3995 13030
rect 4051 13028 4075 13030
rect 4131 13028 4137 13030
rect 3829 13019 4137 13028
rect 3829 11996 4137 12005
rect 3829 11994 3835 11996
rect 3891 11994 3915 11996
rect 3971 11994 3995 11996
rect 4051 11994 4075 11996
rect 4131 11994 4137 11996
rect 3891 11942 3893 11994
rect 4073 11942 4075 11994
rect 3829 11940 3835 11942
rect 3891 11940 3915 11942
rect 3971 11940 3995 11942
rect 4051 11940 4075 11942
rect 4131 11940 4137 11942
rect 3829 11931 4137 11940
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7886 2820 8230
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 3620 6914 3648 10474
rect 3712 7546 3740 11698
rect 3829 10908 4137 10917
rect 3829 10906 3835 10908
rect 3891 10906 3915 10908
rect 3971 10906 3995 10908
rect 4051 10906 4075 10908
rect 4131 10906 4137 10908
rect 3891 10854 3893 10906
rect 4073 10854 4075 10906
rect 3829 10852 3835 10854
rect 3891 10852 3915 10854
rect 3971 10852 3995 10854
rect 4051 10852 4075 10854
rect 4131 10852 4137 10854
rect 3829 10843 4137 10852
rect 4816 10266 4844 13194
rect 5368 12918 5396 16934
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5828 14482 5856 16526
rect 6196 15502 6224 17002
rect 6184 15496 6236 15502
rect 6184 15438 6236 15444
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5828 13462 5856 14418
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5736 11354 5764 13262
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 3829 9820 4137 9829
rect 3829 9818 3835 9820
rect 3891 9818 3915 9820
rect 3971 9818 3995 9820
rect 4051 9818 4075 9820
rect 4131 9818 4137 9820
rect 3891 9766 3893 9818
rect 4073 9766 4075 9818
rect 3829 9764 3835 9766
rect 3891 9764 3915 9766
rect 3971 9764 3995 9766
rect 4051 9764 4075 9766
rect 4131 9764 4137 9766
rect 3829 9755 4137 9764
rect 3829 8732 4137 8741
rect 3829 8730 3835 8732
rect 3891 8730 3915 8732
rect 3971 8730 3995 8732
rect 4051 8730 4075 8732
rect 4131 8730 4137 8732
rect 3891 8678 3893 8730
rect 4073 8678 4075 8730
rect 3829 8676 3835 8678
rect 3891 8676 3915 8678
rect 3971 8676 3995 8678
rect 4051 8676 4075 8678
rect 4131 8676 4137 8678
rect 3829 8667 4137 8676
rect 3829 7644 4137 7653
rect 3829 7642 3835 7644
rect 3891 7642 3915 7644
rect 3971 7642 3995 7644
rect 4051 7642 4075 7644
rect 4131 7642 4137 7644
rect 3891 7590 3893 7642
rect 4073 7590 4075 7642
rect 3829 7588 3835 7590
rect 3891 7588 3915 7590
rect 3971 7588 3995 7590
rect 4051 7588 4075 7590
rect 4131 7588 4137 7590
rect 3829 7579 4137 7588
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3620 6886 3740 6914
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 3712 4690 3740 6886
rect 3829 6556 4137 6565
rect 3829 6554 3835 6556
rect 3891 6554 3915 6556
rect 3971 6554 3995 6556
rect 4051 6554 4075 6556
rect 4131 6554 4137 6556
rect 3891 6502 3893 6554
rect 4073 6502 4075 6554
rect 3829 6500 3835 6502
rect 3891 6500 3915 6502
rect 3971 6500 3995 6502
rect 4051 6500 4075 6502
rect 4131 6500 4137 6502
rect 3829 6491 4137 6500
rect 3829 5468 4137 5477
rect 3829 5466 3835 5468
rect 3891 5466 3915 5468
rect 3971 5466 3995 5468
rect 4051 5466 4075 5468
rect 4131 5466 4137 5468
rect 3891 5414 3893 5466
rect 4073 5414 4075 5466
rect 3829 5412 3835 5414
rect 3891 5412 3915 5414
rect 3971 5412 3995 5414
rect 4051 5412 4075 5414
rect 4131 5412 4137 5414
rect 3829 5403 4137 5412
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 5828 4622 5856 13398
rect 6196 13190 6224 15438
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 8022 6224 13126
rect 6840 9178 6868 17138
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 8036 9586 8064 17274
rect 15016 17264 15068 17270
rect 15016 17206 15068 17212
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 15028 16590 15056 17206
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15120 16658 15148 17138
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15212 16794 15240 16934
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15016 16584 15068 16590
rect 15016 16526 15068 16532
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 8268 16348 8576 16357
rect 8268 16346 8274 16348
rect 8330 16346 8354 16348
rect 8410 16346 8434 16348
rect 8490 16346 8514 16348
rect 8570 16346 8576 16348
rect 8330 16294 8332 16346
rect 8512 16294 8514 16346
rect 8268 16292 8274 16294
rect 8330 16292 8354 16294
rect 8410 16292 8434 16294
rect 8490 16292 8514 16294
rect 8570 16292 8576 16294
rect 8268 16283 8576 16292
rect 8268 15260 8576 15269
rect 8268 15258 8274 15260
rect 8330 15258 8354 15260
rect 8410 15258 8434 15260
rect 8490 15258 8514 15260
rect 8570 15258 8576 15260
rect 8330 15206 8332 15258
rect 8512 15206 8514 15258
rect 8268 15204 8274 15206
rect 8330 15204 8354 15206
rect 8410 15204 8434 15206
rect 8490 15204 8514 15206
rect 8570 15204 8576 15206
rect 8268 15195 8576 15204
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 11354 8156 14282
rect 8268 14172 8576 14181
rect 8268 14170 8274 14172
rect 8330 14170 8354 14172
rect 8410 14170 8434 14172
rect 8490 14170 8514 14172
rect 8570 14170 8576 14172
rect 8330 14118 8332 14170
rect 8512 14118 8514 14170
rect 8268 14116 8274 14118
rect 8330 14116 8354 14118
rect 8410 14116 8434 14118
rect 8490 14116 8514 14118
rect 8570 14116 8576 14118
rect 8268 14107 8576 14116
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8268 13084 8576 13093
rect 8268 13082 8274 13084
rect 8330 13082 8354 13084
rect 8410 13082 8434 13084
rect 8490 13082 8514 13084
rect 8570 13082 8576 13084
rect 8330 13030 8332 13082
rect 8512 13030 8514 13082
rect 8268 13028 8274 13030
rect 8330 13028 8354 13030
rect 8410 13028 8434 13030
rect 8490 13028 8514 13030
rect 8570 13028 8576 13030
rect 8268 13019 8576 13028
rect 8268 11996 8576 12005
rect 8268 11994 8274 11996
rect 8330 11994 8354 11996
rect 8410 11994 8434 11996
rect 8490 11994 8514 11996
rect 8570 11994 8576 11996
rect 8330 11942 8332 11994
rect 8512 11942 8514 11994
rect 8268 11940 8274 11942
rect 8330 11940 8354 11942
rect 8410 11940 8434 11942
rect 8490 11940 8514 11942
rect 8570 11940 8576 11942
rect 8268 11931 8576 11940
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 7484 8430 7512 9454
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 5710 6960 7686
rect 8128 7410 8156 11290
rect 8268 10908 8576 10917
rect 8268 10906 8274 10908
rect 8330 10906 8354 10908
rect 8410 10906 8434 10908
rect 8490 10906 8514 10908
rect 8570 10906 8576 10908
rect 8330 10854 8332 10906
rect 8512 10854 8514 10906
rect 8268 10852 8274 10854
rect 8330 10852 8354 10854
rect 8410 10852 8434 10854
rect 8490 10852 8514 10854
rect 8570 10852 8576 10854
rect 8268 10843 8576 10852
rect 8268 9820 8576 9829
rect 8268 9818 8274 9820
rect 8330 9818 8354 9820
rect 8410 9818 8434 9820
rect 8490 9818 8514 9820
rect 8570 9818 8576 9820
rect 8330 9766 8332 9818
rect 8512 9766 8514 9818
rect 8268 9764 8274 9766
rect 8330 9764 8354 9766
rect 8410 9764 8434 9766
rect 8490 9764 8514 9766
rect 8570 9764 8576 9766
rect 8268 9755 8576 9764
rect 9048 9654 9076 13874
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 11072 9518 11100 16390
rect 12707 16348 13015 16357
rect 12707 16346 12713 16348
rect 12769 16346 12793 16348
rect 12849 16346 12873 16348
rect 12929 16346 12953 16348
rect 13009 16346 13015 16348
rect 12769 16294 12771 16346
rect 12951 16294 12953 16346
rect 12707 16292 12713 16294
rect 12769 16292 12793 16294
rect 12849 16292 12873 16294
rect 12929 16292 12953 16294
rect 13009 16292 13015 16294
rect 12707 16283 13015 16292
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 15028 15434 15056 16526
rect 15212 16114 15240 16730
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15304 15502 15332 16458
rect 17146 16348 17454 16357
rect 17146 16346 17152 16348
rect 17208 16346 17232 16348
rect 17288 16346 17312 16348
rect 17368 16346 17392 16348
rect 17448 16346 17454 16348
rect 17208 16294 17210 16346
rect 17390 16294 17392 16346
rect 17146 16292 17152 16294
rect 17208 16292 17232 16294
rect 17288 16292 17312 16294
rect 17368 16292 17392 16294
rect 17448 16292 17454 16294
rect 17146 16283 17454 16292
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 12707 15260 13015 15269
rect 12707 15258 12713 15260
rect 12769 15258 12793 15260
rect 12849 15258 12873 15260
rect 12929 15258 12953 15260
rect 13009 15258 13015 15260
rect 12769 15206 12771 15258
rect 12951 15206 12953 15258
rect 12707 15204 12713 15206
rect 12769 15204 12793 15206
rect 12849 15204 12873 15206
rect 12929 15204 12953 15206
rect 13009 15204 13015 15206
rect 12707 15195 13015 15204
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 12707 14172 13015 14181
rect 12707 14170 12713 14172
rect 12769 14170 12793 14172
rect 12849 14170 12873 14172
rect 12929 14170 12953 14172
rect 13009 14170 13015 14172
rect 12769 14118 12771 14170
rect 12951 14118 12953 14170
rect 12707 14116 12713 14118
rect 12769 14116 12793 14118
rect 12849 14116 12873 14118
rect 12929 14116 12953 14118
rect 13009 14116 13015 14118
rect 12707 14107 13015 14116
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 12707 13084 13015 13093
rect 12707 13082 12713 13084
rect 12769 13082 12793 13084
rect 12849 13082 12873 13084
rect 12929 13082 12953 13084
rect 13009 13082 13015 13084
rect 12769 13030 12771 13082
rect 12951 13030 12953 13082
rect 12707 13028 12713 13030
rect 12769 13028 12793 13030
rect 12849 13028 12873 13030
rect 12929 13028 12953 13030
rect 13009 13028 13015 13030
rect 12707 13019 13015 13028
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 12707 11996 13015 12005
rect 12707 11994 12713 11996
rect 12769 11994 12793 11996
rect 12849 11994 12873 11996
rect 12929 11994 12953 11996
rect 13009 11994 13015 11996
rect 12769 11942 12771 11994
rect 12951 11942 12953 11994
rect 12707 11940 12713 11942
rect 12769 11940 12793 11942
rect 12849 11940 12873 11942
rect 12929 11940 12953 11942
rect 13009 11940 13015 11942
rect 12707 11931 13015 11940
rect 12047 11452 12355 11461
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 12707 10908 13015 10917
rect 12707 10906 12713 10908
rect 12769 10906 12793 10908
rect 12849 10906 12873 10908
rect 12929 10906 12953 10908
rect 13009 10906 13015 10908
rect 12769 10854 12771 10906
rect 12951 10854 12953 10906
rect 12707 10852 12713 10854
rect 12769 10852 12793 10854
rect 12849 10852 12873 10854
rect 12929 10852 12953 10854
rect 13009 10852 13015 10854
rect 12707 10843 13015 10852
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 12707 9820 13015 9829
rect 12707 9818 12713 9820
rect 12769 9818 12793 9820
rect 12849 9818 12873 9820
rect 12929 9818 12953 9820
rect 13009 9818 13015 9820
rect 12769 9766 12771 9818
rect 12951 9766 12953 9818
rect 12707 9764 12713 9766
rect 12769 9764 12793 9766
rect 12849 9764 12873 9766
rect 12929 9764 12953 9766
rect 13009 9764 13015 9766
rect 12707 9755 13015 9764
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 8268 8732 8576 8741
rect 8268 8730 8274 8732
rect 8330 8730 8354 8732
rect 8410 8730 8434 8732
rect 8490 8730 8514 8732
rect 8570 8730 8576 8732
rect 8330 8678 8332 8730
rect 8512 8678 8514 8730
rect 8268 8676 8274 8678
rect 8330 8676 8354 8678
rect 8410 8676 8434 8678
rect 8490 8676 8514 8678
rect 8570 8676 8576 8678
rect 8268 8667 8576 8676
rect 12707 8732 13015 8741
rect 12707 8730 12713 8732
rect 12769 8730 12793 8732
rect 12849 8730 12873 8732
rect 12929 8730 12953 8732
rect 13009 8730 13015 8732
rect 12769 8678 12771 8730
rect 12951 8678 12953 8730
rect 12707 8676 12713 8678
rect 12769 8676 12793 8678
rect 12849 8676 12873 8678
rect 12929 8676 12953 8678
rect 13009 8676 13015 8678
rect 12707 8667 13015 8676
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 9128 8016 9180 8022
rect 9128 7958 9180 7964
rect 8268 7644 8576 7653
rect 8268 7642 8274 7644
rect 8330 7642 8354 7644
rect 8410 7642 8434 7644
rect 8490 7642 8514 7644
rect 8570 7642 8576 7644
rect 8330 7590 8332 7642
rect 8512 7590 8514 7642
rect 8268 7588 8274 7590
rect 8330 7588 8354 7590
rect 8410 7588 8434 7590
rect 8490 7588 8514 7590
rect 8570 7588 8576 7590
rect 8268 7579 8576 7588
rect 9140 7410 9168 7958
rect 12707 7644 13015 7653
rect 12707 7642 12713 7644
rect 12769 7642 12793 7644
rect 12849 7642 12873 7644
rect 12929 7642 12953 7644
rect 13009 7642 13015 7644
rect 12769 7590 12771 7642
rect 12951 7590 12953 7642
rect 12707 7588 12713 7590
rect 12769 7588 12793 7590
rect 12849 7588 12873 7590
rect 12929 7588 12953 7590
rect 13009 7588 13015 7590
rect 12707 7579 13015 7588
rect 14108 7410 14136 15370
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 8268 6556 8576 6565
rect 8268 6554 8274 6556
rect 8330 6554 8354 6556
rect 8410 6554 8434 6556
rect 8490 6554 8514 6556
rect 8570 6554 8576 6556
rect 8330 6502 8332 6554
rect 8512 6502 8514 6554
rect 8268 6500 8274 6502
rect 8330 6500 8354 6502
rect 8410 6500 8434 6502
rect 8490 6500 8514 6502
rect 8570 6500 8576 6502
rect 8268 6491 8576 6500
rect 12707 6556 13015 6565
rect 12707 6554 12713 6556
rect 12769 6554 12793 6556
rect 12849 6554 12873 6556
rect 12929 6554 12953 6556
rect 13009 6554 13015 6556
rect 12769 6502 12771 6554
rect 12951 6502 12953 6554
rect 12707 6500 12713 6502
rect 12769 6500 12793 6502
rect 12849 6500 12873 6502
rect 12929 6500 12953 6502
rect 13009 6500 13015 6502
rect 12707 6491 13015 6500
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 8268 5468 8576 5477
rect 8268 5466 8274 5468
rect 8330 5466 8354 5468
rect 8410 5466 8434 5468
rect 8490 5466 8514 5468
rect 8570 5466 8576 5468
rect 8330 5414 8332 5466
rect 8512 5414 8514 5466
rect 8268 5412 8274 5414
rect 8330 5412 8354 5414
rect 8410 5412 8434 5414
rect 8490 5412 8514 5414
rect 8570 5412 8576 5414
rect 8268 5403 8576 5412
rect 12707 5468 13015 5477
rect 12707 5466 12713 5468
rect 12769 5466 12793 5468
rect 12849 5466 12873 5468
rect 12929 5466 12953 5468
rect 13009 5466 13015 5468
rect 12769 5414 12771 5466
rect 12951 5414 12953 5466
rect 12707 5412 12713 5414
rect 12769 5412 12793 5414
rect 12849 5412 12873 5414
rect 12929 5412 12953 5414
rect 13009 5412 13015 5414
rect 12707 5403 13015 5412
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 13832 4486 13860 5646
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 3829 4380 4137 4389
rect 3829 4378 3835 4380
rect 3891 4378 3915 4380
rect 3971 4378 3995 4380
rect 4051 4378 4075 4380
rect 4131 4378 4137 4380
rect 3891 4326 3893 4378
rect 4073 4326 4075 4378
rect 3829 4324 3835 4326
rect 3891 4324 3915 4326
rect 3971 4324 3995 4326
rect 4051 4324 4075 4326
rect 4131 4324 4137 4326
rect 3829 4315 4137 4324
rect 8268 4380 8576 4389
rect 8268 4378 8274 4380
rect 8330 4378 8354 4380
rect 8410 4378 8434 4380
rect 8490 4378 8514 4380
rect 8570 4378 8576 4380
rect 8330 4326 8332 4378
rect 8512 4326 8514 4378
rect 8268 4324 8274 4326
rect 8330 4324 8354 4326
rect 8410 4324 8434 4326
rect 8490 4324 8514 4326
rect 8570 4324 8576 4326
rect 8268 4315 8576 4324
rect 12707 4380 13015 4389
rect 12707 4378 12713 4380
rect 12769 4378 12793 4380
rect 12849 4378 12873 4380
rect 12929 4378 12953 4380
rect 13009 4378 13015 4380
rect 12769 4326 12771 4378
rect 12951 4326 12953 4378
rect 12707 4324 12713 4326
rect 12769 4324 12793 4326
rect 12849 4324 12873 4326
rect 12929 4324 12953 4326
rect 13009 4324 13015 4326
rect 12707 4315 13015 4324
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 3829 3292 4137 3301
rect 3829 3290 3835 3292
rect 3891 3290 3915 3292
rect 3971 3290 3995 3292
rect 4051 3290 4075 3292
rect 4131 3290 4137 3292
rect 3891 3238 3893 3290
rect 4073 3238 4075 3290
rect 3829 3236 3835 3238
rect 3891 3236 3915 3238
rect 3971 3236 3995 3238
rect 4051 3236 4075 3238
rect 4131 3236 4137 3238
rect 3829 3227 4137 3236
rect 8268 3292 8576 3301
rect 8268 3290 8274 3292
rect 8330 3290 8354 3292
rect 8410 3290 8434 3292
rect 8490 3290 8514 3292
rect 8570 3290 8576 3292
rect 8330 3238 8332 3290
rect 8512 3238 8514 3290
rect 8268 3236 8274 3238
rect 8330 3236 8354 3238
rect 8410 3236 8434 3238
rect 8490 3236 8514 3238
rect 8570 3236 8576 3238
rect 8268 3227 8576 3236
rect 12707 3292 13015 3301
rect 12707 3290 12713 3292
rect 12769 3290 12793 3292
rect 12849 3290 12873 3292
rect 12929 3290 12953 3292
rect 13009 3290 13015 3292
rect 12769 3238 12771 3290
rect 12951 3238 12953 3290
rect 12707 3236 12713 3238
rect 12769 3236 12793 3238
rect 12849 3236 12873 3238
rect 12929 3236 12953 3238
rect 13009 3236 13015 3238
rect 12707 3227 13015 3236
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 13924 2446 13952 7210
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 15396 2378 15424 15302
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 16960 13258 16988 14350
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 17052 7274 17080 15982
rect 17146 15260 17454 15269
rect 17146 15258 17152 15260
rect 17208 15258 17232 15260
rect 17288 15258 17312 15260
rect 17368 15258 17392 15260
rect 17448 15258 17454 15260
rect 17208 15206 17210 15258
rect 17390 15206 17392 15258
rect 17146 15204 17152 15206
rect 17208 15204 17232 15206
rect 17288 15204 17312 15206
rect 17368 15204 17392 15206
rect 17448 15204 17454 15206
rect 17146 15195 17454 15204
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 17146 14172 17454 14181
rect 17146 14170 17152 14172
rect 17208 14170 17232 14172
rect 17288 14170 17312 14172
rect 17368 14170 17392 14172
rect 17448 14170 17454 14172
rect 17208 14118 17210 14170
rect 17390 14118 17392 14170
rect 17146 14116 17152 14118
rect 17208 14116 17232 14118
rect 17288 14116 17312 14118
rect 17368 14116 17392 14118
rect 17448 14116 17454 14118
rect 17146 14107 17454 14116
rect 18156 13938 18184 14418
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18420 14272 18472 14278
rect 18420 14214 18472 14220
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17146 13084 17454 13093
rect 17146 13082 17152 13084
rect 17208 13082 17232 13084
rect 17288 13082 17312 13084
rect 17368 13082 17392 13084
rect 17448 13082 17454 13084
rect 17208 13030 17210 13082
rect 17390 13030 17392 13082
rect 17146 13028 17152 13030
rect 17208 13028 17232 13030
rect 17288 13028 17312 13030
rect 17368 13028 17392 13030
rect 17448 13028 17454 13030
rect 17146 13019 17454 13028
rect 17146 11996 17454 12005
rect 17146 11994 17152 11996
rect 17208 11994 17232 11996
rect 17288 11994 17312 11996
rect 17368 11994 17392 11996
rect 17448 11994 17454 11996
rect 17208 11942 17210 11994
rect 17390 11942 17392 11994
rect 17146 11940 17152 11942
rect 17208 11940 17232 11942
rect 17288 11940 17312 11942
rect 17368 11940 17392 11942
rect 17448 11940 17454 11942
rect 17146 11931 17454 11940
rect 17146 10908 17454 10917
rect 17146 10906 17152 10908
rect 17208 10906 17232 10908
rect 17288 10906 17312 10908
rect 17368 10906 17392 10908
rect 17448 10906 17454 10908
rect 17208 10854 17210 10906
rect 17390 10854 17392 10906
rect 17146 10852 17152 10854
rect 17208 10852 17232 10854
rect 17288 10852 17312 10854
rect 17368 10852 17392 10854
rect 17448 10852 17454 10854
rect 17146 10843 17454 10852
rect 17146 9820 17454 9829
rect 17146 9818 17152 9820
rect 17208 9818 17232 9820
rect 17288 9818 17312 9820
rect 17368 9818 17392 9820
rect 17448 9818 17454 9820
rect 17208 9766 17210 9818
rect 17390 9766 17392 9818
rect 17146 9764 17152 9766
rect 17208 9764 17232 9766
rect 17288 9764 17312 9766
rect 17368 9764 17392 9766
rect 17448 9764 17454 9766
rect 17146 9755 17454 9764
rect 17146 8732 17454 8741
rect 17146 8730 17152 8732
rect 17208 8730 17232 8732
rect 17288 8730 17312 8732
rect 17368 8730 17392 8732
rect 17448 8730 17454 8732
rect 17208 8678 17210 8730
rect 17390 8678 17392 8730
rect 17146 8676 17152 8678
rect 17208 8676 17232 8678
rect 17288 8676 17312 8678
rect 17368 8676 17392 8678
rect 17448 8676 17454 8678
rect 17146 8667 17454 8676
rect 17146 7644 17454 7653
rect 17146 7642 17152 7644
rect 17208 7642 17232 7644
rect 17288 7642 17312 7644
rect 17368 7642 17392 7644
rect 17448 7642 17454 7644
rect 17208 7590 17210 7642
rect 17390 7590 17392 7642
rect 17146 7588 17152 7590
rect 17208 7588 17232 7590
rect 17288 7588 17312 7590
rect 17368 7588 17392 7590
rect 17448 7588 17454 7590
rect 17146 7579 17454 7588
rect 17512 7342 17540 13806
rect 18432 7818 18460 14214
rect 18524 13938 18552 14350
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18524 13394 18552 13874
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17040 7268 17092 7274
rect 17040 7210 17092 7216
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 17146 6556 17454 6565
rect 17146 6554 17152 6556
rect 17208 6554 17232 6556
rect 17288 6554 17312 6556
rect 17368 6554 17392 6556
rect 17448 6554 17454 6556
rect 17208 6502 17210 6554
rect 17390 6502 17392 6554
rect 17146 6500 17152 6502
rect 17208 6500 17232 6502
rect 17288 6500 17312 6502
rect 17368 6500 17392 6502
rect 17448 6500 17454 6502
rect 17146 6491 17454 6500
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 17512 5710 17540 7278
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17146 5468 17454 5477
rect 17146 5466 17152 5468
rect 17208 5466 17232 5468
rect 17288 5466 17312 5468
rect 17368 5466 17392 5468
rect 17448 5466 17454 5468
rect 17208 5414 17210 5466
rect 17390 5414 17392 5466
rect 17146 5412 17152 5414
rect 17208 5412 17232 5414
rect 17288 5412 17312 5414
rect 17368 5412 17392 5414
rect 17448 5412 17454 5414
rect 17146 5403 17454 5412
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 17146 4380 17454 4389
rect 17146 4378 17152 4380
rect 17208 4378 17232 4380
rect 17288 4378 17312 4380
rect 17368 4378 17392 4380
rect 17448 4378 17454 4380
rect 17208 4326 17210 4378
rect 17390 4326 17392 4378
rect 17146 4324 17152 4326
rect 17208 4324 17232 4326
rect 17288 4324 17312 4326
rect 17368 4324 17392 4326
rect 17448 4324 17454 4326
rect 17146 4315 17454 4324
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 17146 3292 17454 3301
rect 17146 3290 17152 3292
rect 17208 3290 17232 3292
rect 17288 3290 17312 3292
rect 17368 3290 17392 3292
rect 17448 3290 17454 3292
rect 17208 3238 17210 3290
rect 17390 3238 17392 3290
rect 17146 3236 17152 3238
rect 17208 3236 17232 3238
rect 17288 3236 17312 3238
rect 17368 3236 17392 3238
rect 17448 3236 17454 3238
rect 17146 3227 17454 3236
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 15384 2372 15436 2378
rect 15384 2314 15436 2320
rect 3829 2204 4137 2213
rect 3829 2202 3835 2204
rect 3891 2202 3915 2204
rect 3971 2202 3995 2204
rect 4051 2202 4075 2204
rect 4131 2202 4137 2204
rect 3891 2150 3893 2202
rect 4073 2150 4075 2202
rect 3829 2148 3835 2150
rect 3891 2148 3915 2150
rect 3971 2148 3995 2150
rect 4051 2148 4075 2150
rect 4131 2148 4137 2150
rect 3829 2139 4137 2148
rect 8268 2204 8576 2213
rect 8268 2202 8274 2204
rect 8330 2202 8354 2204
rect 8410 2202 8434 2204
rect 8490 2202 8514 2204
rect 8570 2202 8576 2204
rect 8330 2150 8332 2202
rect 8512 2150 8514 2202
rect 8268 2148 8274 2150
rect 8330 2148 8354 2150
rect 8410 2148 8434 2150
rect 8490 2148 8514 2150
rect 8570 2148 8576 2150
rect 8268 2139 8576 2148
rect 12707 2204 13015 2213
rect 12707 2202 12713 2204
rect 12769 2202 12793 2204
rect 12849 2202 12873 2204
rect 12929 2202 12953 2204
rect 13009 2202 13015 2204
rect 12769 2150 12771 2202
rect 12951 2150 12953 2202
rect 12707 2148 12713 2150
rect 12769 2148 12793 2150
rect 12849 2148 12873 2150
rect 12929 2148 12953 2150
rect 13009 2148 13015 2150
rect 12707 2139 13015 2148
rect 17146 2204 17454 2213
rect 17146 2202 17152 2204
rect 17208 2202 17232 2204
rect 17288 2202 17312 2204
rect 17368 2202 17392 2204
rect 17448 2202 17454 2204
rect 17208 2150 17210 2202
rect 17390 2150 17392 2202
rect 17146 2148 17152 2150
rect 17208 2148 17232 2150
rect 17288 2148 17312 2150
rect 17368 2148 17392 2150
rect 17448 2148 17454 2150
rect 17146 2139 17454 2148
<< via2 >>
rect 3835 17434 3891 17436
rect 3915 17434 3971 17436
rect 3995 17434 4051 17436
rect 4075 17434 4131 17436
rect 3835 17382 3881 17434
rect 3881 17382 3891 17434
rect 3915 17382 3945 17434
rect 3945 17382 3957 17434
rect 3957 17382 3971 17434
rect 3995 17382 4009 17434
rect 4009 17382 4021 17434
rect 4021 17382 4051 17434
rect 4075 17382 4085 17434
rect 4085 17382 4131 17434
rect 3835 17380 3891 17382
rect 3915 17380 3971 17382
rect 3995 17380 4051 17382
rect 4075 17380 4131 17382
rect 8274 17434 8330 17436
rect 8354 17434 8410 17436
rect 8434 17434 8490 17436
rect 8514 17434 8570 17436
rect 8274 17382 8320 17434
rect 8320 17382 8330 17434
rect 8354 17382 8384 17434
rect 8384 17382 8396 17434
rect 8396 17382 8410 17434
rect 8434 17382 8448 17434
rect 8448 17382 8460 17434
rect 8460 17382 8490 17434
rect 8514 17382 8524 17434
rect 8524 17382 8570 17434
rect 8274 17380 8330 17382
rect 8354 17380 8410 17382
rect 8434 17380 8490 17382
rect 8514 17380 8570 17382
rect 12713 17434 12769 17436
rect 12793 17434 12849 17436
rect 12873 17434 12929 17436
rect 12953 17434 13009 17436
rect 12713 17382 12759 17434
rect 12759 17382 12769 17434
rect 12793 17382 12823 17434
rect 12823 17382 12835 17434
rect 12835 17382 12849 17434
rect 12873 17382 12887 17434
rect 12887 17382 12899 17434
rect 12899 17382 12929 17434
rect 12953 17382 12963 17434
rect 12963 17382 13009 17434
rect 12713 17380 12769 17382
rect 12793 17380 12849 17382
rect 12873 17380 12929 17382
rect 12953 17380 13009 17382
rect 17152 17434 17208 17436
rect 17232 17434 17288 17436
rect 17312 17434 17368 17436
rect 17392 17434 17448 17436
rect 17152 17382 17198 17434
rect 17198 17382 17208 17434
rect 17232 17382 17262 17434
rect 17262 17382 17274 17434
rect 17274 17382 17288 17434
rect 17312 17382 17326 17434
rect 17326 17382 17338 17434
rect 17338 17382 17368 17434
rect 17392 17382 17402 17434
rect 17402 17382 17448 17434
rect 17152 17380 17208 17382
rect 17232 17380 17288 17382
rect 17312 17380 17368 17382
rect 17392 17380 17448 17382
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 1490 15000 1546 15056
rect 846 14492 848 14512
rect 848 14492 900 14512
rect 900 14492 902 14512
rect 846 14456 902 14492
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 846 13132 848 13152
rect 848 13132 900 13152
rect 900 13132 902 13152
rect 846 13096 902 13132
rect 1490 12280 1546 12336
rect 846 11464 902 11520
rect 1490 10920 1546 10976
rect 846 10376 902 10432
rect 1398 9560 1454 9616
rect 846 9016 902 9072
rect 1398 8200 1454 8256
rect 846 7692 848 7712
rect 848 7692 900 7712
rect 900 7692 902 7712
rect 846 7656 902 7692
rect 1490 6840 1546 6896
rect 846 6296 902 6352
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 846 4936 902 4992
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 3835 16346 3891 16348
rect 3915 16346 3971 16348
rect 3995 16346 4051 16348
rect 4075 16346 4131 16348
rect 3835 16294 3881 16346
rect 3881 16294 3891 16346
rect 3915 16294 3945 16346
rect 3945 16294 3957 16346
rect 3957 16294 3971 16346
rect 3995 16294 4009 16346
rect 4009 16294 4021 16346
rect 4021 16294 4051 16346
rect 4075 16294 4085 16346
rect 4085 16294 4131 16346
rect 3835 16292 3891 16294
rect 3915 16292 3971 16294
rect 3995 16292 4051 16294
rect 4075 16292 4131 16294
rect 3835 15258 3891 15260
rect 3915 15258 3971 15260
rect 3995 15258 4051 15260
rect 4075 15258 4131 15260
rect 3835 15206 3881 15258
rect 3881 15206 3891 15258
rect 3915 15206 3945 15258
rect 3945 15206 3957 15258
rect 3957 15206 3971 15258
rect 3995 15206 4009 15258
rect 4009 15206 4021 15258
rect 4021 15206 4051 15258
rect 4075 15206 4085 15258
rect 4085 15206 4131 15258
rect 3835 15204 3891 15206
rect 3915 15204 3971 15206
rect 3995 15204 4051 15206
rect 4075 15204 4131 15206
rect 3835 14170 3891 14172
rect 3915 14170 3971 14172
rect 3995 14170 4051 14172
rect 4075 14170 4131 14172
rect 3835 14118 3881 14170
rect 3881 14118 3891 14170
rect 3915 14118 3945 14170
rect 3945 14118 3957 14170
rect 3957 14118 3971 14170
rect 3995 14118 4009 14170
rect 4009 14118 4021 14170
rect 4021 14118 4051 14170
rect 4075 14118 4085 14170
rect 4085 14118 4131 14170
rect 3835 14116 3891 14118
rect 3915 14116 3971 14118
rect 3995 14116 4051 14118
rect 4075 14116 4131 14118
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 3835 13082 3891 13084
rect 3915 13082 3971 13084
rect 3995 13082 4051 13084
rect 4075 13082 4131 13084
rect 3835 13030 3881 13082
rect 3881 13030 3891 13082
rect 3915 13030 3945 13082
rect 3945 13030 3957 13082
rect 3957 13030 3971 13082
rect 3995 13030 4009 13082
rect 4009 13030 4021 13082
rect 4021 13030 4051 13082
rect 4075 13030 4085 13082
rect 4085 13030 4131 13082
rect 3835 13028 3891 13030
rect 3915 13028 3971 13030
rect 3995 13028 4051 13030
rect 4075 13028 4131 13030
rect 3835 11994 3891 11996
rect 3915 11994 3971 11996
rect 3995 11994 4051 11996
rect 4075 11994 4131 11996
rect 3835 11942 3881 11994
rect 3881 11942 3891 11994
rect 3915 11942 3945 11994
rect 3945 11942 3957 11994
rect 3957 11942 3971 11994
rect 3995 11942 4009 11994
rect 4009 11942 4021 11994
rect 4021 11942 4051 11994
rect 4075 11942 4085 11994
rect 4085 11942 4131 11994
rect 3835 11940 3891 11942
rect 3915 11940 3971 11942
rect 3995 11940 4051 11942
rect 4075 11940 4131 11942
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 3835 10906 3891 10908
rect 3915 10906 3971 10908
rect 3995 10906 4051 10908
rect 4075 10906 4131 10908
rect 3835 10854 3881 10906
rect 3881 10854 3891 10906
rect 3915 10854 3945 10906
rect 3945 10854 3957 10906
rect 3957 10854 3971 10906
rect 3995 10854 4009 10906
rect 4009 10854 4021 10906
rect 4021 10854 4051 10906
rect 4075 10854 4085 10906
rect 4085 10854 4131 10906
rect 3835 10852 3891 10854
rect 3915 10852 3971 10854
rect 3995 10852 4051 10854
rect 4075 10852 4131 10854
rect 3835 9818 3891 9820
rect 3915 9818 3971 9820
rect 3995 9818 4051 9820
rect 4075 9818 4131 9820
rect 3835 9766 3881 9818
rect 3881 9766 3891 9818
rect 3915 9766 3945 9818
rect 3945 9766 3957 9818
rect 3957 9766 3971 9818
rect 3995 9766 4009 9818
rect 4009 9766 4021 9818
rect 4021 9766 4051 9818
rect 4075 9766 4085 9818
rect 4085 9766 4131 9818
rect 3835 9764 3891 9766
rect 3915 9764 3971 9766
rect 3995 9764 4051 9766
rect 4075 9764 4131 9766
rect 3835 8730 3891 8732
rect 3915 8730 3971 8732
rect 3995 8730 4051 8732
rect 4075 8730 4131 8732
rect 3835 8678 3881 8730
rect 3881 8678 3891 8730
rect 3915 8678 3945 8730
rect 3945 8678 3957 8730
rect 3957 8678 3971 8730
rect 3995 8678 4009 8730
rect 4009 8678 4021 8730
rect 4021 8678 4051 8730
rect 4075 8678 4085 8730
rect 4085 8678 4131 8730
rect 3835 8676 3891 8678
rect 3915 8676 3971 8678
rect 3995 8676 4051 8678
rect 4075 8676 4131 8678
rect 3835 7642 3891 7644
rect 3915 7642 3971 7644
rect 3995 7642 4051 7644
rect 4075 7642 4131 7644
rect 3835 7590 3881 7642
rect 3881 7590 3891 7642
rect 3915 7590 3945 7642
rect 3945 7590 3957 7642
rect 3957 7590 3971 7642
rect 3995 7590 4009 7642
rect 4009 7590 4021 7642
rect 4021 7590 4051 7642
rect 4075 7590 4085 7642
rect 4085 7590 4131 7642
rect 3835 7588 3891 7590
rect 3915 7588 3971 7590
rect 3995 7588 4051 7590
rect 4075 7588 4131 7590
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 3835 6554 3891 6556
rect 3915 6554 3971 6556
rect 3995 6554 4051 6556
rect 4075 6554 4131 6556
rect 3835 6502 3881 6554
rect 3881 6502 3891 6554
rect 3915 6502 3945 6554
rect 3945 6502 3957 6554
rect 3957 6502 3971 6554
rect 3995 6502 4009 6554
rect 4009 6502 4021 6554
rect 4021 6502 4051 6554
rect 4075 6502 4085 6554
rect 4085 6502 4131 6554
rect 3835 6500 3891 6502
rect 3915 6500 3971 6502
rect 3995 6500 4051 6502
rect 4075 6500 4131 6502
rect 3835 5466 3891 5468
rect 3915 5466 3971 5468
rect 3995 5466 4051 5468
rect 4075 5466 4131 5468
rect 3835 5414 3881 5466
rect 3881 5414 3891 5466
rect 3915 5414 3945 5466
rect 3945 5414 3957 5466
rect 3957 5414 3971 5466
rect 3995 5414 4009 5466
rect 4009 5414 4021 5466
rect 4021 5414 4051 5466
rect 4075 5414 4085 5466
rect 4085 5414 4131 5466
rect 3835 5412 3891 5414
rect 3915 5412 3971 5414
rect 3995 5412 4051 5414
rect 4075 5412 4131 5414
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 8274 16346 8330 16348
rect 8354 16346 8410 16348
rect 8434 16346 8490 16348
rect 8514 16346 8570 16348
rect 8274 16294 8320 16346
rect 8320 16294 8330 16346
rect 8354 16294 8384 16346
rect 8384 16294 8396 16346
rect 8396 16294 8410 16346
rect 8434 16294 8448 16346
rect 8448 16294 8460 16346
rect 8460 16294 8490 16346
rect 8514 16294 8524 16346
rect 8524 16294 8570 16346
rect 8274 16292 8330 16294
rect 8354 16292 8410 16294
rect 8434 16292 8490 16294
rect 8514 16292 8570 16294
rect 8274 15258 8330 15260
rect 8354 15258 8410 15260
rect 8434 15258 8490 15260
rect 8514 15258 8570 15260
rect 8274 15206 8320 15258
rect 8320 15206 8330 15258
rect 8354 15206 8384 15258
rect 8384 15206 8396 15258
rect 8396 15206 8410 15258
rect 8434 15206 8448 15258
rect 8448 15206 8460 15258
rect 8460 15206 8490 15258
rect 8514 15206 8524 15258
rect 8524 15206 8570 15258
rect 8274 15204 8330 15206
rect 8354 15204 8410 15206
rect 8434 15204 8490 15206
rect 8514 15204 8570 15206
rect 8274 14170 8330 14172
rect 8354 14170 8410 14172
rect 8434 14170 8490 14172
rect 8514 14170 8570 14172
rect 8274 14118 8320 14170
rect 8320 14118 8330 14170
rect 8354 14118 8384 14170
rect 8384 14118 8396 14170
rect 8396 14118 8410 14170
rect 8434 14118 8448 14170
rect 8448 14118 8460 14170
rect 8460 14118 8490 14170
rect 8514 14118 8524 14170
rect 8524 14118 8570 14170
rect 8274 14116 8330 14118
rect 8354 14116 8410 14118
rect 8434 14116 8490 14118
rect 8514 14116 8570 14118
rect 8274 13082 8330 13084
rect 8354 13082 8410 13084
rect 8434 13082 8490 13084
rect 8514 13082 8570 13084
rect 8274 13030 8320 13082
rect 8320 13030 8330 13082
rect 8354 13030 8384 13082
rect 8384 13030 8396 13082
rect 8396 13030 8410 13082
rect 8434 13030 8448 13082
rect 8448 13030 8460 13082
rect 8460 13030 8490 13082
rect 8514 13030 8524 13082
rect 8524 13030 8570 13082
rect 8274 13028 8330 13030
rect 8354 13028 8410 13030
rect 8434 13028 8490 13030
rect 8514 13028 8570 13030
rect 8274 11994 8330 11996
rect 8354 11994 8410 11996
rect 8434 11994 8490 11996
rect 8514 11994 8570 11996
rect 8274 11942 8320 11994
rect 8320 11942 8330 11994
rect 8354 11942 8384 11994
rect 8384 11942 8396 11994
rect 8396 11942 8410 11994
rect 8434 11942 8448 11994
rect 8448 11942 8460 11994
rect 8460 11942 8490 11994
rect 8514 11942 8524 11994
rect 8524 11942 8570 11994
rect 8274 11940 8330 11942
rect 8354 11940 8410 11942
rect 8434 11940 8490 11942
rect 8514 11940 8570 11942
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 8274 10906 8330 10908
rect 8354 10906 8410 10908
rect 8434 10906 8490 10908
rect 8514 10906 8570 10908
rect 8274 10854 8320 10906
rect 8320 10854 8330 10906
rect 8354 10854 8384 10906
rect 8384 10854 8396 10906
rect 8396 10854 8410 10906
rect 8434 10854 8448 10906
rect 8448 10854 8460 10906
rect 8460 10854 8490 10906
rect 8514 10854 8524 10906
rect 8524 10854 8570 10906
rect 8274 10852 8330 10854
rect 8354 10852 8410 10854
rect 8434 10852 8490 10854
rect 8514 10852 8570 10854
rect 8274 9818 8330 9820
rect 8354 9818 8410 9820
rect 8434 9818 8490 9820
rect 8514 9818 8570 9820
rect 8274 9766 8320 9818
rect 8320 9766 8330 9818
rect 8354 9766 8384 9818
rect 8384 9766 8396 9818
rect 8396 9766 8410 9818
rect 8434 9766 8448 9818
rect 8448 9766 8460 9818
rect 8460 9766 8490 9818
rect 8514 9766 8524 9818
rect 8524 9766 8570 9818
rect 8274 9764 8330 9766
rect 8354 9764 8410 9766
rect 8434 9764 8490 9766
rect 8514 9764 8570 9766
rect 12713 16346 12769 16348
rect 12793 16346 12849 16348
rect 12873 16346 12929 16348
rect 12953 16346 13009 16348
rect 12713 16294 12759 16346
rect 12759 16294 12769 16346
rect 12793 16294 12823 16346
rect 12823 16294 12835 16346
rect 12835 16294 12849 16346
rect 12873 16294 12887 16346
rect 12887 16294 12899 16346
rect 12899 16294 12929 16346
rect 12953 16294 12963 16346
rect 12963 16294 13009 16346
rect 12713 16292 12769 16294
rect 12793 16292 12849 16294
rect 12873 16292 12929 16294
rect 12953 16292 13009 16294
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 17152 16346 17208 16348
rect 17232 16346 17288 16348
rect 17312 16346 17368 16348
rect 17392 16346 17448 16348
rect 17152 16294 17198 16346
rect 17198 16294 17208 16346
rect 17232 16294 17262 16346
rect 17262 16294 17274 16346
rect 17274 16294 17288 16346
rect 17312 16294 17326 16346
rect 17326 16294 17338 16346
rect 17338 16294 17368 16346
rect 17392 16294 17402 16346
rect 17402 16294 17448 16346
rect 17152 16292 17208 16294
rect 17232 16292 17288 16294
rect 17312 16292 17368 16294
rect 17392 16292 17448 16294
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 12713 15258 12769 15260
rect 12793 15258 12849 15260
rect 12873 15258 12929 15260
rect 12953 15258 13009 15260
rect 12713 15206 12759 15258
rect 12759 15206 12769 15258
rect 12793 15206 12823 15258
rect 12823 15206 12835 15258
rect 12835 15206 12849 15258
rect 12873 15206 12887 15258
rect 12887 15206 12899 15258
rect 12899 15206 12929 15258
rect 12953 15206 12963 15258
rect 12963 15206 13009 15258
rect 12713 15204 12769 15206
rect 12793 15204 12849 15206
rect 12873 15204 12929 15206
rect 12953 15204 13009 15206
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 12713 14170 12769 14172
rect 12793 14170 12849 14172
rect 12873 14170 12929 14172
rect 12953 14170 13009 14172
rect 12713 14118 12759 14170
rect 12759 14118 12769 14170
rect 12793 14118 12823 14170
rect 12823 14118 12835 14170
rect 12835 14118 12849 14170
rect 12873 14118 12887 14170
rect 12887 14118 12899 14170
rect 12899 14118 12929 14170
rect 12953 14118 12963 14170
rect 12963 14118 13009 14170
rect 12713 14116 12769 14118
rect 12793 14116 12849 14118
rect 12873 14116 12929 14118
rect 12953 14116 13009 14118
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 12713 13082 12769 13084
rect 12793 13082 12849 13084
rect 12873 13082 12929 13084
rect 12953 13082 13009 13084
rect 12713 13030 12759 13082
rect 12759 13030 12769 13082
rect 12793 13030 12823 13082
rect 12823 13030 12835 13082
rect 12835 13030 12849 13082
rect 12873 13030 12887 13082
rect 12887 13030 12899 13082
rect 12899 13030 12929 13082
rect 12953 13030 12963 13082
rect 12963 13030 13009 13082
rect 12713 13028 12769 13030
rect 12793 13028 12849 13030
rect 12873 13028 12929 13030
rect 12953 13028 13009 13030
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 12713 11994 12769 11996
rect 12793 11994 12849 11996
rect 12873 11994 12929 11996
rect 12953 11994 13009 11996
rect 12713 11942 12759 11994
rect 12759 11942 12769 11994
rect 12793 11942 12823 11994
rect 12823 11942 12835 11994
rect 12835 11942 12849 11994
rect 12873 11942 12887 11994
rect 12887 11942 12899 11994
rect 12899 11942 12929 11994
rect 12953 11942 12963 11994
rect 12963 11942 13009 11994
rect 12713 11940 12769 11942
rect 12793 11940 12849 11942
rect 12873 11940 12929 11942
rect 12953 11940 13009 11942
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 12713 10906 12769 10908
rect 12793 10906 12849 10908
rect 12873 10906 12929 10908
rect 12953 10906 13009 10908
rect 12713 10854 12759 10906
rect 12759 10854 12769 10906
rect 12793 10854 12823 10906
rect 12823 10854 12835 10906
rect 12835 10854 12849 10906
rect 12873 10854 12887 10906
rect 12887 10854 12899 10906
rect 12899 10854 12929 10906
rect 12953 10854 12963 10906
rect 12963 10854 13009 10906
rect 12713 10852 12769 10854
rect 12793 10852 12849 10854
rect 12873 10852 12929 10854
rect 12953 10852 13009 10854
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 12713 9818 12769 9820
rect 12793 9818 12849 9820
rect 12873 9818 12929 9820
rect 12953 9818 13009 9820
rect 12713 9766 12759 9818
rect 12759 9766 12769 9818
rect 12793 9766 12823 9818
rect 12823 9766 12835 9818
rect 12835 9766 12849 9818
rect 12873 9766 12887 9818
rect 12887 9766 12899 9818
rect 12899 9766 12929 9818
rect 12953 9766 12963 9818
rect 12963 9766 13009 9818
rect 12713 9764 12769 9766
rect 12793 9764 12849 9766
rect 12873 9764 12929 9766
rect 12953 9764 13009 9766
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 8274 8730 8330 8732
rect 8354 8730 8410 8732
rect 8434 8730 8490 8732
rect 8514 8730 8570 8732
rect 8274 8678 8320 8730
rect 8320 8678 8330 8730
rect 8354 8678 8384 8730
rect 8384 8678 8396 8730
rect 8396 8678 8410 8730
rect 8434 8678 8448 8730
rect 8448 8678 8460 8730
rect 8460 8678 8490 8730
rect 8514 8678 8524 8730
rect 8524 8678 8570 8730
rect 8274 8676 8330 8678
rect 8354 8676 8410 8678
rect 8434 8676 8490 8678
rect 8514 8676 8570 8678
rect 12713 8730 12769 8732
rect 12793 8730 12849 8732
rect 12873 8730 12929 8732
rect 12953 8730 13009 8732
rect 12713 8678 12759 8730
rect 12759 8678 12769 8730
rect 12793 8678 12823 8730
rect 12823 8678 12835 8730
rect 12835 8678 12849 8730
rect 12873 8678 12887 8730
rect 12887 8678 12899 8730
rect 12899 8678 12929 8730
rect 12953 8678 12963 8730
rect 12963 8678 13009 8730
rect 12713 8676 12769 8678
rect 12793 8676 12849 8678
rect 12873 8676 12929 8678
rect 12953 8676 13009 8678
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 8274 7642 8330 7644
rect 8354 7642 8410 7644
rect 8434 7642 8490 7644
rect 8514 7642 8570 7644
rect 8274 7590 8320 7642
rect 8320 7590 8330 7642
rect 8354 7590 8384 7642
rect 8384 7590 8396 7642
rect 8396 7590 8410 7642
rect 8434 7590 8448 7642
rect 8448 7590 8460 7642
rect 8460 7590 8490 7642
rect 8514 7590 8524 7642
rect 8524 7590 8570 7642
rect 8274 7588 8330 7590
rect 8354 7588 8410 7590
rect 8434 7588 8490 7590
rect 8514 7588 8570 7590
rect 12713 7642 12769 7644
rect 12793 7642 12849 7644
rect 12873 7642 12929 7644
rect 12953 7642 13009 7644
rect 12713 7590 12759 7642
rect 12759 7590 12769 7642
rect 12793 7590 12823 7642
rect 12823 7590 12835 7642
rect 12835 7590 12849 7642
rect 12873 7590 12887 7642
rect 12887 7590 12899 7642
rect 12899 7590 12929 7642
rect 12953 7590 12963 7642
rect 12963 7590 13009 7642
rect 12713 7588 12769 7590
rect 12793 7588 12849 7590
rect 12873 7588 12929 7590
rect 12953 7588 13009 7590
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 8274 6554 8330 6556
rect 8354 6554 8410 6556
rect 8434 6554 8490 6556
rect 8514 6554 8570 6556
rect 8274 6502 8320 6554
rect 8320 6502 8330 6554
rect 8354 6502 8384 6554
rect 8384 6502 8396 6554
rect 8396 6502 8410 6554
rect 8434 6502 8448 6554
rect 8448 6502 8460 6554
rect 8460 6502 8490 6554
rect 8514 6502 8524 6554
rect 8524 6502 8570 6554
rect 8274 6500 8330 6502
rect 8354 6500 8410 6502
rect 8434 6500 8490 6502
rect 8514 6500 8570 6502
rect 12713 6554 12769 6556
rect 12793 6554 12849 6556
rect 12873 6554 12929 6556
rect 12953 6554 13009 6556
rect 12713 6502 12759 6554
rect 12759 6502 12769 6554
rect 12793 6502 12823 6554
rect 12823 6502 12835 6554
rect 12835 6502 12849 6554
rect 12873 6502 12887 6554
rect 12887 6502 12899 6554
rect 12899 6502 12929 6554
rect 12953 6502 12963 6554
rect 12963 6502 13009 6554
rect 12713 6500 12769 6502
rect 12793 6500 12849 6502
rect 12873 6500 12929 6502
rect 12953 6500 13009 6502
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 8274 5466 8330 5468
rect 8354 5466 8410 5468
rect 8434 5466 8490 5468
rect 8514 5466 8570 5468
rect 8274 5414 8320 5466
rect 8320 5414 8330 5466
rect 8354 5414 8384 5466
rect 8384 5414 8396 5466
rect 8396 5414 8410 5466
rect 8434 5414 8448 5466
rect 8448 5414 8460 5466
rect 8460 5414 8490 5466
rect 8514 5414 8524 5466
rect 8524 5414 8570 5466
rect 8274 5412 8330 5414
rect 8354 5412 8410 5414
rect 8434 5412 8490 5414
rect 8514 5412 8570 5414
rect 12713 5466 12769 5468
rect 12793 5466 12849 5468
rect 12873 5466 12929 5468
rect 12953 5466 13009 5468
rect 12713 5414 12759 5466
rect 12759 5414 12769 5466
rect 12793 5414 12823 5466
rect 12823 5414 12835 5466
rect 12835 5414 12849 5466
rect 12873 5414 12887 5466
rect 12887 5414 12899 5466
rect 12899 5414 12929 5466
rect 12953 5414 12963 5466
rect 12963 5414 13009 5466
rect 12713 5412 12769 5414
rect 12793 5412 12849 5414
rect 12873 5412 12929 5414
rect 12953 5412 13009 5414
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 3835 4378 3891 4380
rect 3915 4378 3971 4380
rect 3995 4378 4051 4380
rect 4075 4378 4131 4380
rect 3835 4326 3881 4378
rect 3881 4326 3891 4378
rect 3915 4326 3945 4378
rect 3945 4326 3957 4378
rect 3957 4326 3971 4378
rect 3995 4326 4009 4378
rect 4009 4326 4021 4378
rect 4021 4326 4051 4378
rect 4075 4326 4085 4378
rect 4085 4326 4131 4378
rect 3835 4324 3891 4326
rect 3915 4324 3971 4326
rect 3995 4324 4051 4326
rect 4075 4324 4131 4326
rect 8274 4378 8330 4380
rect 8354 4378 8410 4380
rect 8434 4378 8490 4380
rect 8514 4378 8570 4380
rect 8274 4326 8320 4378
rect 8320 4326 8330 4378
rect 8354 4326 8384 4378
rect 8384 4326 8396 4378
rect 8396 4326 8410 4378
rect 8434 4326 8448 4378
rect 8448 4326 8460 4378
rect 8460 4326 8490 4378
rect 8514 4326 8524 4378
rect 8524 4326 8570 4378
rect 8274 4324 8330 4326
rect 8354 4324 8410 4326
rect 8434 4324 8490 4326
rect 8514 4324 8570 4326
rect 12713 4378 12769 4380
rect 12793 4378 12849 4380
rect 12873 4378 12929 4380
rect 12953 4378 13009 4380
rect 12713 4326 12759 4378
rect 12759 4326 12769 4378
rect 12793 4326 12823 4378
rect 12823 4326 12835 4378
rect 12835 4326 12849 4378
rect 12873 4326 12887 4378
rect 12887 4326 12899 4378
rect 12899 4326 12929 4378
rect 12953 4326 12963 4378
rect 12963 4326 13009 4378
rect 12713 4324 12769 4326
rect 12793 4324 12849 4326
rect 12873 4324 12929 4326
rect 12953 4324 13009 4326
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 3835 3290 3891 3292
rect 3915 3290 3971 3292
rect 3995 3290 4051 3292
rect 4075 3290 4131 3292
rect 3835 3238 3881 3290
rect 3881 3238 3891 3290
rect 3915 3238 3945 3290
rect 3945 3238 3957 3290
rect 3957 3238 3971 3290
rect 3995 3238 4009 3290
rect 4009 3238 4021 3290
rect 4021 3238 4051 3290
rect 4075 3238 4085 3290
rect 4085 3238 4131 3290
rect 3835 3236 3891 3238
rect 3915 3236 3971 3238
rect 3995 3236 4051 3238
rect 4075 3236 4131 3238
rect 8274 3290 8330 3292
rect 8354 3290 8410 3292
rect 8434 3290 8490 3292
rect 8514 3290 8570 3292
rect 8274 3238 8320 3290
rect 8320 3238 8330 3290
rect 8354 3238 8384 3290
rect 8384 3238 8396 3290
rect 8396 3238 8410 3290
rect 8434 3238 8448 3290
rect 8448 3238 8460 3290
rect 8460 3238 8490 3290
rect 8514 3238 8524 3290
rect 8524 3238 8570 3290
rect 8274 3236 8330 3238
rect 8354 3236 8410 3238
rect 8434 3236 8490 3238
rect 8514 3236 8570 3238
rect 12713 3290 12769 3292
rect 12793 3290 12849 3292
rect 12873 3290 12929 3292
rect 12953 3290 13009 3292
rect 12713 3238 12759 3290
rect 12759 3238 12769 3290
rect 12793 3238 12823 3290
rect 12823 3238 12835 3290
rect 12835 3238 12849 3290
rect 12873 3238 12887 3290
rect 12887 3238 12899 3290
rect 12899 3238 12929 3290
rect 12953 3238 12963 3290
rect 12963 3238 13009 3290
rect 12713 3236 12769 3238
rect 12793 3236 12849 3238
rect 12873 3236 12929 3238
rect 12953 3236 13009 3238
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 17152 15258 17208 15260
rect 17232 15258 17288 15260
rect 17312 15258 17368 15260
rect 17392 15258 17448 15260
rect 17152 15206 17198 15258
rect 17198 15206 17208 15258
rect 17232 15206 17262 15258
rect 17262 15206 17274 15258
rect 17274 15206 17288 15258
rect 17312 15206 17326 15258
rect 17326 15206 17338 15258
rect 17338 15206 17368 15258
rect 17392 15206 17402 15258
rect 17402 15206 17448 15258
rect 17152 15204 17208 15206
rect 17232 15204 17288 15206
rect 17312 15204 17368 15206
rect 17392 15204 17448 15206
rect 17152 14170 17208 14172
rect 17232 14170 17288 14172
rect 17312 14170 17368 14172
rect 17392 14170 17448 14172
rect 17152 14118 17198 14170
rect 17198 14118 17208 14170
rect 17232 14118 17262 14170
rect 17262 14118 17274 14170
rect 17274 14118 17288 14170
rect 17312 14118 17326 14170
rect 17326 14118 17338 14170
rect 17338 14118 17368 14170
rect 17392 14118 17402 14170
rect 17402 14118 17448 14170
rect 17152 14116 17208 14118
rect 17232 14116 17288 14118
rect 17312 14116 17368 14118
rect 17392 14116 17448 14118
rect 17152 13082 17208 13084
rect 17232 13082 17288 13084
rect 17312 13082 17368 13084
rect 17392 13082 17448 13084
rect 17152 13030 17198 13082
rect 17198 13030 17208 13082
rect 17232 13030 17262 13082
rect 17262 13030 17274 13082
rect 17274 13030 17288 13082
rect 17312 13030 17326 13082
rect 17326 13030 17338 13082
rect 17338 13030 17368 13082
rect 17392 13030 17402 13082
rect 17402 13030 17448 13082
rect 17152 13028 17208 13030
rect 17232 13028 17288 13030
rect 17312 13028 17368 13030
rect 17392 13028 17448 13030
rect 17152 11994 17208 11996
rect 17232 11994 17288 11996
rect 17312 11994 17368 11996
rect 17392 11994 17448 11996
rect 17152 11942 17198 11994
rect 17198 11942 17208 11994
rect 17232 11942 17262 11994
rect 17262 11942 17274 11994
rect 17274 11942 17288 11994
rect 17312 11942 17326 11994
rect 17326 11942 17338 11994
rect 17338 11942 17368 11994
rect 17392 11942 17402 11994
rect 17402 11942 17448 11994
rect 17152 11940 17208 11942
rect 17232 11940 17288 11942
rect 17312 11940 17368 11942
rect 17392 11940 17448 11942
rect 17152 10906 17208 10908
rect 17232 10906 17288 10908
rect 17312 10906 17368 10908
rect 17392 10906 17448 10908
rect 17152 10854 17198 10906
rect 17198 10854 17208 10906
rect 17232 10854 17262 10906
rect 17262 10854 17274 10906
rect 17274 10854 17288 10906
rect 17312 10854 17326 10906
rect 17326 10854 17338 10906
rect 17338 10854 17368 10906
rect 17392 10854 17402 10906
rect 17402 10854 17448 10906
rect 17152 10852 17208 10854
rect 17232 10852 17288 10854
rect 17312 10852 17368 10854
rect 17392 10852 17448 10854
rect 17152 9818 17208 9820
rect 17232 9818 17288 9820
rect 17312 9818 17368 9820
rect 17392 9818 17448 9820
rect 17152 9766 17198 9818
rect 17198 9766 17208 9818
rect 17232 9766 17262 9818
rect 17262 9766 17274 9818
rect 17274 9766 17288 9818
rect 17312 9766 17326 9818
rect 17326 9766 17338 9818
rect 17338 9766 17368 9818
rect 17392 9766 17402 9818
rect 17402 9766 17448 9818
rect 17152 9764 17208 9766
rect 17232 9764 17288 9766
rect 17312 9764 17368 9766
rect 17392 9764 17448 9766
rect 17152 8730 17208 8732
rect 17232 8730 17288 8732
rect 17312 8730 17368 8732
rect 17392 8730 17448 8732
rect 17152 8678 17198 8730
rect 17198 8678 17208 8730
rect 17232 8678 17262 8730
rect 17262 8678 17274 8730
rect 17274 8678 17288 8730
rect 17312 8678 17326 8730
rect 17326 8678 17338 8730
rect 17338 8678 17368 8730
rect 17392 8678 17402 8730
rect 17402 8678 17448 8730
rect 17152 8676 17208 8678
rect 17232 8676 17288 8678
rect 17312 8676 17368 8678
rect 17392 8676 17448 8678
rect 17152 7642 17208 7644
rect 17232 7642 17288 7644
rect 17312 7642 17368 7644
rect 17392 7642 17448 7644
rect 17152 7590 17198 7642
rect 17198 7590 17208 7642
rect 17232 7590 17262 7642
rect 17262 7590 17274 7642
rect 17274 7590 17288 7642
rect 17312 7590 17326 7642
rect 17326 7590 17338 7642
rect 17338 7590 17368 7642
rect 17392 7590 17402 7642
rect 17402 7590 17448 7642
rect 17152 7588 17208 7590
rect 17232 7588 17288 7590
rect 17312 7588 17368 7590
rect 17392 7588 17448 7590
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 17152 6554 17208 6556
rect 17232 6554 17288 6556
rect 17312 6554 17368 6556
rect 17392 6554 17448 6556
rect 17152 6502 17198 6554
rect 17198 6502 17208 6554
rect 17232 6502 17262 6554
rect 17262 6502 17274 6554
rect 17274 6502 17288 6554
rect 17312 6502 17326 6554
rect 17326 6502 17338 6554
rect 17338 6502 17368 6554
rect 17392 6502 17402 6554
rect 17402 6502 17448 6554
rect 17152 6500 17208 6502
rect 17232 6500 17288 6502
rect 17312 6500 17368 6502
rect 17392 6500 17448 6502
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 17152 5466 17208 5468
rect 17232 5466 17288 5468
rect 17312 5466 17368 5468
rect 17392 5466 17448 5468
rect 17152 5414 17198 5466
rect 17198 5414 17208 5466
rect 17232 5414 17262 5466
rect 17262 5414 17274 5466
rect 17274 5414 17288 5466
rect 17312 5414 17326 5466
rect 17326 5414 17338 5466
rect 17338 5414 17368 5466
rect 17392 5414 17402 5466
rect 17402 5414 17448 5466
rect 17152 5412 17208 5414
rect 17232 5412 17288 5414
rect 17312 5412 17368 5414
rect 17392 5412 17448 5414
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 17152 4378 17208 4380
rect 17232 4378 17288 4380
rect 17312 4378 17368 4380
rect 17392 4378 17448 4380
rect 17152 4326 17198 4378
rect 17198 4326 17208 4378
rect 17232 4326 17262 4378
rect 17262 4326 17274 4378
rect 17274 4326 17288 4378
rect 17312 4326 17326 4378
rect 17326 4326 17338 4378
rect 17338 4326 17368 4378
rect 17392 4326 17402 4378
rect 17402 4326 17448 4378
rect 17152 4324 17208 4326
rect 17232 4324 17288 4326
rect 17312 4324 17368 4326
rect 17392 4324 17448 4326
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 17152 3290 17208 3292
rect 17232 3290 17288 3292
rect 17312 3290 17368 3292
rect 17392 3290 17448 3292
rect 17152 3238 17198 3290
rect 17198 3238 17208 3290
rect 17232 3238 17262 3290
rect 17262 3238 17274 3290
rect 17274 3238 17288 3290
rect 17312 3238 17326 3290
rect 17326 3238 17338 3290
rect 17338 3238 17368 3290
rect 17392 3238 17402 3290
rect 17402 3238 17448 3290
rect 17152 3236 17208 3238
rect 17232 3236 17288 3238
rect 17312 3236 17368 3238
rect 17392 3236 17448 3238
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 3835 2202 3891 2204
rect 3915 2202 3971 2204
rect 3995 2202 4051 2204
rect 4075 2202 4131 2204
rect 3835 2150 3881 2202
rect 3881 2150 3891 2202
rect 3915 2150 3945 2202
rect 3945 2150 3957 2202
rect 3957 2150 3971 2202
rect 3995 2150 4009 2202
rect 4009 2150 4021 2202
rect 4021 2150 4051 2202
rect 4075 2150 4085 2202
rect 4085 2150 4131 2202
rect 3835 2148 3891 2150
rect 3915 2148 3971 2150
rect 3995 2148 4051 2150
rect 4075 2148 4131 2150
rect 8274 2202 8330 2204
rect 8354 2202 8410 2204
rect 8434 2202 8490 2204
rect 8514 2202 8570 2204
rect 8274 2150 8320 2202
rect 8320 2150 8330 2202
rect 8354 2150 8384 2202
rect 8384 2150 8396 2202
rect 8396 2150 8410 2202
rect 8434 2150 8448 2202
rect 8448 2150 8460 2202
rect 8460 2150 8490 2202
rect 8514 2150 8524 2202
rect 8524 2150 8570 2202
rect 8274 2148 8330 2150
rect 8354 2148 8410 2150
rect 8434 2148 8490 2150
rect 8514 2148 8570 2150
rect 12713 2202 12769 2204
rect 12793 2202 12849 2204
rect 12873 2202 12929 2204
rect 12953 2202 13009 2204
rect 12713 2150 12759 2202
rect 12759 2150 12769 2202
rect 12793 2150 12823 2202
rect 12823 2150 12835 2202
rect 12835 2150 12849 2202
rect 12873 2150 12887 2202
rect 12887 2150 12899 2202
rect 12899 2150 12929 2202
rect 12953 2150 12963 2202
rect 12963 2150 13009 2202
rect 12713 2148 12769 2150
rect 12793 2148 12849 2150
rect 12873 2148 12929 2150
rect 12953 2148 13009 2150
rect 17152 2202 17208 2204
rect 17232 2202 17288 2204
rect 17312 2202 17368 2204
rect 17392 2202 17448 2204
rect 17152 2150 17198 2202
rect 17198 2150 17208 2202
rect 17232 2150 17262 2202
rect 17262 2150 17274 2202
rect 17274 2150 17288 2202
rect 17312 2150 17326 2202
rect 17326 2150 17338 2202
rect 17338 2150 17368 2202
rect 17392 2150 17402 2202
rect 17402 2150 17448 2202
rect 17152 2148 17208 2150
rect 17232 2148 17288 2150
rect 17312 2148 17368 2150
rect 17392 2148 17448 2150
<< metal3 >>
rect 3825 17440 4141 17441
rect 3825 17376 3831 17440
rect 3895 17376 3911 17440
rect 3975 17376 3991 17440
rect 4055 17376 4071 17440
rect 4135 17376 4141 17440
rect 3825 17375 4141 17376
rect 8264 17440 8580 17441
rect 8264 17376 8270 17440
rect 8334 17376 8350 17440
rect 8414 17376 8430 17440
rect 8494 17376 8510 17440
rect 8574 17376 8580 17440
rect 8264 17375 8580 17376
rect 12703 17440 13019 17441
rect 12703 17376 12709 17440
rect 12773 17376 12789 17440
rect 12853 17376 12869 17440
rect 12933 17376 12949 17440
rect 13013 17376 13019 17440
rect 12703 17375 13019 17376
rect 17142 17440 17458 17441
rect 17142 17376 17148 17440
rect 17212 17376 17228 17440
rect 17292 17376 17308 17440
rect 17372 17376 17388 17440
rect 17452 17376 17458 17440
rect 17142 17375 17458 17376
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 16482 16831 16798 16832
rect 3825 16352 4141 16353
rect 3825 16288 3831 16352
rect 3895 16288 3911 16352
rect 3975 16288 3991 16352
rect 4055 16288 4071 16352
rect 4135 16288 4141 16352
rect 3825 16287 4141 16288
rect 8264 16352 8580 16353
rect 8264 16288 8270 16352
rect 8334 16288 8350 16352
rect 8414 16288 8430 16352
rect 8494 16288 8510 16352
rect 8574 16288 8580 16352
rect 8264 16287 8580 16288
rect 12703 16352 13019 16353
rect 12703 16288 12709 16352
rect 12773 16288 12789 16352
rect 12853 16288 12869 16352
rect 12933 16288 12949 16352
rect 13013 16288 13019 16352
rect 12703 16287 13019 16288
rect 17142 16352 17458 16353
rect 17142 16288 17148 16352
rect 17212 16288 17228 16352
rect 17292 16288 17308 16352
rect 17372 16288 17388 16352
rect 17452 16288 17458 16352
rect 17142 16287 17458 16288
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 3825 15264 4141 15265
rect 3825 15200 3831 15264
rect 3895 15200 3911 15264
rect 3975 15200 3991 15264
rect 4055 15200 4071 15264
rect 4135 15200 4141 15264
rect 3825 15199 4141 15200
rect 8264 15264 8580 15265
rect 8264 15200 8270 15264
rect 8334 15200 8350 15264
rect 8414 15200 8430 15264
rect 8494 15200 8510 15264
rect 8574 15200 8580 15264
rect 8264 15199 8580 15200
rect 12703 15264 13019 15265
rect 12703 15200 12709 15264
rect 12773 15200 12789 15264
rect 12853 15200 12869 15264
rect 12933 15200 12949 15264
rect 13013 15200 13019 15264
rect 12703 15199 13019 15200
rect 17142 15264 17458 15265
rect 17142 15200 17148 15264
rect 17212 15200 17228 15264
rect 17292 15200 17308 15264
rect 17372 15200 17388 15264
rect 17452 15200 17458 15264
rect 17142 15199 17458 15200
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 3165 14720 3481 14721
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 0 14288 800 14318
rect 3825 14176 4141 14177
rect 3825 14112 3831 14176
rect 3895 14112 3911 14176
rect 3975 14112 3991 14176
rect 4055 14112 4071 14176
rect 4135 14112 4141 14176
rect 3825 14111 4141 14112
rect 8264 14176 8580 14177
rect 8264 14112 8270 14176
rect 8334 14112 8350 14176
rect 8414 14112 8430 14176
rect 8494 14112 8510 14176
rect 8574 14112 8580 14176
rect 8264 14111 8580 14112
rect 12703 14176 13019 14177
rect 12703 14112 12709 14176
rect 12773 14112 12789 14176
rect 12853 14112 12869 14176
rect 12933 14112 12949 14176
rect 13013 14112 13019 14176
rect 12703 14111 13019 14112
rect 17142 14176 17458 14177
rect 17142 14112 17148 14176
rect 17212 14112 17228 14176
rect 17292 14112 17308 14176
rect 17372 14112 17388 14176
rect 17452 14112 17458 14176
rect 17142 14111 17458 14112
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 3825 13088 4141 13089
rect 3825 13024 3831 13088
rect 3895 13024 3911 13088
rect 3975 13024 3991 13088
rect 4055 13024 4071 13088
rect 4135 13024 4141 13088
rect 3825 13023 4141 13024
rect 8264 13088 8580 13089
rect 8264 13024 8270 13088
rect 8334 13024 8350 13088
rect 8414 13024 8430 13088
rect 8494 13024 8510 13088
rect 8574 13024 8580 13088
rect 8264 13023 8580 13024
rect 12703 13088 13019 13089
rect 12703 13024 12709 13088
rect 12773 13024 12789 13088
rect 12853 13024 12869 13088
rect 12933 13024 12949 13088
rect 13013 13024 13019 13088
rect 12703 13023 13019 13024
rect 17142 13088 17458 13089
rect 17142 13024 17148 13088
rect 17212 13024 17228 13088
rect 17292 13024 17308 13088
rect 17372 13024 17388 13088
rect 17452 13024 17458 13088
rect 17142 13023 17458 13024
rect 0 12928 800 12958
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 3825 12000 4141 12001
rect 3825 11936 3831 12000
rect 3895 11936 3911 12000
rect 3975 11936 3991 12000
rect 4055 11936 4071 12000
rect 4135 11936 4141 12000
rect 3825 11935 4141 11936
rect 8264 12000 8580 12001
rect 8264 11936 8270 12000
rect 8334 11936 8350 12000
rect 8414 11936 8430 12000
rect 8494 11936 8510 12000
rect 8574 11936 8580 12000
rect 8264 11935 8580 11936
rect 12703 12000 13019 12001
rect 12703 11936 12709 12000
rect 12773 11936 12789 12000
rect 12853 11936 12869 12000
rect 12933 11936 12949 12000
rect 13013 11936 13019 12000
rect 12703 11935 13019 11936
rect 17142 12000 17458 12001
rect 17142 11936 17148 12000
rect 17212 11936 17228 12000
rect 17292 11936 17308 12000
rect 17372 11936 17388 12000
rect 17452 11936 17458 12000
rect 17142 11935 17458 11936
rect 0 11658 800 11688
rect 0 11568 858 11658
rect 798 11525 858 11568
rect 798 11520 907 11525
rect 798 11464 846 11520
rect 902 11464 907 11520
rect 798 11462 907 11464
rect 841 11459 907 11462
rect 3165 11456 3481 11457
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 3825 10912 4141 10913
rect 3825 10848 3831 10912
rect 3895 10848 3911 10912
rect 3975 10848 3991 10912
rect 4055 10848 4071 10912
rect 4135 10848 4141 10912
rect 3825 10847 4141 10848
rect 8264 10912 8580 10913
rect 8264 10848 8270 10912
rect 8334 10848 8350 10912
rect 8414 10848 8430 10912
rect 8494 10848 8510 10912
rect 8574 10848 8580 10912
rect 8264 10847 8580 10848
rect 12703 10912 13019 10913
rect 12703 10848 12709 10912
rect 12773 10848 12789 10912
rect 12853 10848 12869 10912
rect 12933 10848 12949 10912
rect 13013 10848 13019 10912
rect 12703 10847 13019 10848
rect 17142 10912 17458 10913
rect 17142 10848 17148 10912
rect 17212 10848 17228 10912
rect 17292 10848 17308 10912
rect 17372 10848 17388 10912
rect 17452 10848 17458 10912
rect 17142 10847 17458 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 16482 10303 16798 10304
rect 0 10208 800 10238
rect 3825 9824 4141 9825
rect 3825 9760 3831 9824
rect 3895 9760 3911 9824
rect 3975 9760 3991 9824
rect 4055 9760 4071 9824
rect 4135 9760 4141 9824
rect 3825 9759 4141 9760
rect 8264 9824 8580 9825
rect 8264 9760 8270 9824
rect 8334 9760 8350 9824
rect 8414 9760 8430 9824
rect 8494 9760 8510 9824
rect 8574 9760 8580 9824
rect 8264 9759 8580 9760
rect 12703 9824 13019 9825
rect 12703 9760 12709 9824
rect 12773 9760 12789 9824
rect 12853 9760 12869 9824
rect 12933 9760 12949 9824
rect 13013 9760 13019 9824
rect 12703 9759 13019 9760
rect 17142 9824 17458 9825
rect 17142 9760 17148 9824
rect 17212 9760 17228 9824
rect 17292 9760 17308 9824
rect 17372 9760 17388 9824
rect 17452 9760 17458 9824
rect 17142 9759 17458 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 16482 9215 16798 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 0 8848 800 8878
rect 3825 8736 4141 8737
rect 3825 8672 3831 8736
rect 3895 8672 3911 8736
rect 3975 8672 3991 8736
rect 4055 8672 4071 8736
rect 4135 8672 4141 8736
rect 3825 8671 4141 8672
rect 8264 8736 8580 8737
rect 8264 8672 8270 8736
rect 8334 8672 8350 8736
rect 8414 8672 8430 8736
rect 8494 8672 8510 8736
rect 8574 8672 8580 8736
rect 8264 8671 8580 8672
rect 12703 8736 13019 8737
rect 12703 8672 12709 8736
rect 12773 8672 12789 8736
rect 12853 8672 12869 8736
rect 12933 8672 12949 8736
rect 13013 8672 13019 8736
rect 12703 8671 13019 8672
rect 17142 8736 17458 8737
rect 17142 8672 17148 8736
rect 17212 8672 17228 8736
rect 17292 8672 17308 8736
rect 17372 8672 17388 8736
rect 17452 8672 17458 8736
rect 17142 8671 17458 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 3165 8192 3481 8193
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 3825 7648 4141 7649
rect 3825 7584 3831 7648
rect 3895 7584 3911 7648
rect 3975 7584 3991 7648
rect 4055 7584 4071 7648
rect 4135 7584 4141 7648
rect 3825 7583 4141 7584
rect 8264 7648 8580 7649
rect 8264 7584 8270 7648
rect 8334 7584 8350 7648
rect 8414 7584 8430 7648
rect 8494 7584 8510 7648
rect 8574 7584 8580 7648
rect 8264 7583 8580 7584
rect 12703 7648 13019 7649
rect 12703 7584 12709 7648
rect 12773 7584 12789 7648
rect 12853 7584 12869 7648
rect 12933 7584 12949 7648
rect 13013 7584 13019 7648
rect 12703 7583 13019 7584
rect 17142 7648 17458 7649
rect 17142 7584 17148 7648
rect 17212 7584 17228 7648
rect 17292 7584 17308 7648
rect 17372 7584 17388 7648
rect 17452 7584 17458 7648
rect 17142 7583 17458 7584
rect 0 7488 800 7518
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 3825 6560 4141 6561
rect 3825 6496 3831 6560
rect 3895 6496 3911 6560
rect 3975 6496 3991 6560
rect 4055 6496 4071 6560
rect 4135 6496 4141 6560
rect 3825 6495 4141 6496
rect 8264 6560 8580 6561
rect 8264 6496 8270 6560
rect 8334 6496 8350 6560
rect 8414 6496 8430 6560
rect 8494 6496 8510 6560
rect 8574 6496 8580 6560
rect 8264 6495 8580 6496
rect 12703 6560 13019 6561
rect 12703 6496 12709 6560
rect 12773 6496 12789 6560
rect 12853 6496 12869 6560
rect 12933 6496 12949 6560
rect 13013 6496 13019 6560
rect 12703 6495 13019 6496
rect 17142 6560 17458 6561
rect 17142 6496 17148 6560
rect 17212 6496 17228 6560
rect 17292 6496 17308 6560
rect 17372 6496 17388 6560
rect 17452 6496 17458 6560
rect 17142 6495 17458 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 0 6128 800 6158
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 3825 5472 4141 5473
rect 3825 5408 3831 5472
rect 3895 5408 3911 5472
rect 3975 5408 3991 5472
rect 4055 5408 4071 5472
rect 4135 5408 4141 5472
rect 3825 5407 4141 5408
rect 8264 5472 8580 5473
rect 8264 5408 8270 5472
rect 8334 5408 8350 5472
rect 8414 5408 8430 5472
rect 8494 5408 8510 5472
rect 8574 5408 8580 5472
rect 8264 5407 8580 5408
rect 12703 5472 13019 5473
rect 12703 5408 12709 5472
rect 12773 5408 12789 5472
rect 12853 5408 12869 5472
rect 12933 5408 12949 5472
rect 13013 5408 13019 5472
rect 12703 5407 13019 5408
rect 17142 5472 17458 5473
rect 17142 5408 17148 5472
rect 17212 5408 17228 5472
rect 17292 5408 17308 5472
rect 17372 5408 17388 5472
rect 17452 5408 17458 5472
rect 17142 5407 17458 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 0 4768 800 4798
rect 3825 4384 4141 4385
rect 3825 4320 3831 4384
rect 3895 4320 3911 4384
rect 3975 4320 3991 4384
rect 4055 4320 4071 4384
rect 4135 4320 4141 4384
rect 3825 4319 4141 4320
rect 8264 4384 8580 4385
rect 8264 4320 8270 4384
rect 8334 4320 8350 4384
rect 8414 4320 8430 4384
rect 8494 4320 8510 4384
rect 8574 4320 8580 4384
rect 8264 4319 8580 4320
rect 12703 4384 13019 4385
rect 12703 4320 12709 4384
rect 12773 4320 12789 4384
rect 12853 4320 12869 4384
rect 12933 4320 12949 4384
rect 13013 4320 13019 4384
rect 12703 4319 13019 4320
rect 17142 4384 17458 4385
rect 17142 4320 17148 4384
rect 17212 4320 17228 4384
rect 17292 4320 17308 4384
rect 17372 4320 17388 4384
rect 17452 4320 17458 4384
rect 17142 4319 17458 4320
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 3825 3296 4141 3297
rect 3825 3232 3831 3296
rect 3895 3232 3911 3296
rect 3975 3232 3991 3296
rect 4055 3232 4071 3296
rect 4135 3232 4141 3296
rect 3825 3231 4141 3232
rect 8264 3296 8580 3297
rect 8264 3232 8270 3296
rect 8334 3232 8350 3296
rect 8414 3232 8430 3296
rect 8494 3232 8510 3296
rect 8574 3232 8580 3296
rect 8264 3231 8580 3232
rect 12703 3296 13019 3297
rect 12703 3232 12709 3296
rect 12773 3232 12789 3296
rect 12853 3232 12869 3296
rect 12933 3232 12949 3296
rect 13013 3232 13019 3296
rect 12703 3231 13019 3232
rect 17142 3296 17458 3297
rect 17142 3232 17148 3296
rect 17212 3232 17228 3296
rect 17292 3232 17308 3296
rect 17372 3232 17388 3296
rect 17452 3232 17458 3296
rect 17142 3231 17458 3232
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 3825 2208 4141 2209
rect 3825 2144 3831 2208
rect 3895 2144 3911 2208
rect 3975 2144 3991 2208
rect 4055 2144 4071 2208
rect 4135 2144 4141 2208
rect 3825 2143 4141 2144
rect 8264 2208 8580 2209
rect 8264 2144 8270 2208
rect 8334 2144 8350 2208
rect 8414 2144 8430 2208
rect 8494 2144 8510 2208
rect 8574 2144 8580 2208
rect 8264 2143 8580 2144
rect 12703 2208 13019 2209
rect 12703 2144 12709 2208
rect 12773 2144 12789 2208
rect 12853 2144 12869 2208
rect 12933 2144 12949 2208
rect 13013 2144 13019 2208
rect 12703 2143 13019 2144
rect 17142 2208 17458 2209
rect 17142 2144 17148 2208
rect 17212 2144 17228 2208
rect 17292 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17458 2208
rect 17142 2143 17458 2144
<< via3 >>
rect 3831 17436 3895 17440
rect 3831 17380 3835 17436
rect 3835 17380 3891 17436
rect 3891 17380 3895 17436
rect 3831 17376 3895 17380
rect 3911 17436 3975 17440
rect 3911 17380 3915 17436
rect 3915 17380 3971 17436
rect 3971 17380 3975 17436
rect 3911 17376 3975 17380
rect 3991 17436 4055 17440
rect 3991 17380 3995 17436
rect 3995 17380 4051 17436
rect 4051 17380 4055 17436
rect 3991 17376 4055 17380
rect 4071 17436 4135 17440
rect 4071 17380 4075 17436
rect 4075 17380 4131 17436
rect 4131 17380 4135 17436
rect 4071 17376 4135 17380
rect 8270 17436 8334 17440
rect 8270 17380 8274 17436
rect 8274 17380 8330 17436
rect 8330 17380 8334 17436
rect 8270 17376 8334 17380
rect 8350 17436 8414 17440
rect 8350 17380 8354 17436
rect 8354 17380 8410 17436
rect 8410 17380 8414 17436
rect 8350 17376 8414 17380
rect 8430 17436 8494 17440
rect 8430 17380 8434 17436
rect 8434 17380 8490 17436
rect 8490 17380 8494 17436
rect 8430 17376 8494 17380
rect 8510 17436 8574 17440
rect 8510 17380 8514 17436
rect 8514 17380 8570 17436
rect 8570 17380 8574 17436
rect 8510 17376 8574 17380
rect 12709 17436 12773 17440
rect 12709 17380 12713 17436
rect 12713 17380 12769 17436
rect 12769 17380 12773 17436
rect 12709 17376 12773 17380
rect 12789 17436 12853 17440
rect 12789 17380 12793 17436
rect 12793 17380 12849 17436
rect 12849 17380 12853 17436
rect 12789 17376 12853 17380
rect 12869 17436 12933 17440
rect 12869 17380 12873 17436
rect 12873 17380 12929 17436
rect 12929 17380 12933 17436
rect 12869 17376 12933 17380
rect 12949 17436 13013 17440
rect 12949 17380 12953 17436
rect 12953 17380 13009 17436
rect 13009 17380 13013 17436
rect 12949 17376 13013 17380
rect 17148 17436 17212 17440
rect 17148 17380 17152 17436
rect 17152 17380 17208 17436
rect 17208 17380 17212 17436
rect 17148 17376 17212 17380
rect 17228 17436 17292 17440
rect 17228 17380 17232 17436
rect 17232 17380 17288 17436
rect 17288 17380 17292 17436
rect 17228 17376 17292 17380
rect 17308 17436 17372 17440
rect 17308 17380 17312 17436
rect 17312 17380 17368 17436
rect 17368 17380 17372 17436
rect 17308 17376 17372 17380
rect 17388 17436 17452 17440
rect 17388 17380 17392 17436
rect 17392 17380 17448 17436
rect 17448 17380 17452 17436
rect 17388 17376 17452 17380
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 3831 16348 3895 16352
rect 3831 16292 3835 16348
rect 3835 16292 3891 16348
rect 3891 16292 3895 16348
rect 3831 16288 3895 16292
rect 3911 16348 3975 16352
rect 3911 16292 3915 16348
rect 3915 16292 3971 16348
rect 3971 16292 3975 16348
rect 3911 16288 3975 16292
rect 3991 16348 4055 16352
rect 3991 16292 3995 16348
rect 3995 16292 4051 16348
rect 4051 16292 4055 16348
rect 3991 16288 4055 16292
rect 4071 16348 4135 16352
rect 4071 16292 4075 16348
rect 4075 16292 4131 16348
rect 4131 16292 4135 16348
rect 4071 16288 4135 16292
rect 8270 16348 8334 16352
rect 8270 16292 8274 16348
rect 8274 16292 8330 16348
rect 8330 16292 8334 16348
rect 8270 16288 8334 16292
rect 8350 16348 8414 16352
rect 8350 16292 8354 16348
rect 8354 16292 8410 16348
rect 8410 16292 8414 16348
rect 8350 16288 8414 16292
rect 8430 16348 8494 16352
rect 8430 16292 8434 16348
rect 8434 16292 8490 16348
rect 8490 16292 8494 16348
rect 8430 16288 8494 16292
rect 8510 16348 8574 16352
rect 8510 16292 8514 16348
rect 8514 16292 8570 16348
rect 8570 16292 8574 16348
rect 8510 16288 8574 16292
rect 12709 16348 12773 16352
rect 12709 16292 12713 16348
rect 12713 16292 12769 16348
rect 12769 16292 12773 16348
rect 12709 16288 12773 16292
rect 12789 16348 12853 16352
rect 12789 16292 12793 16348
rect 12793 16292 12849 16348
rect 12849 16292 12853 16348
rect 12789 16288 12853 16292
rect 12869 16348 12933 16352
rect 12869 16292 12873 16348
rect 12873 16292 12929 16348
rect 12929 16292 12933 16348
rect 12869 16288 12933 16292
rect 12949 16348 13013 16352
rect 12949 16292 12953 16348
rect 12953 16292 13009 16348
rect 13009 16292 13013 16348
rect 12949 16288 13013 16292
rect 17148 16348 17212 16352
rect 17148 16292 17152 16348
rect 17152 16292 17208 16348
rect 17208 16292 17212 16348
rect 17148 16288 17212 16292
rect 17228 16348 17292 16352
rect 17228 16292 17232 16348
rect 17232 16292 17288 16348
rect 17288 16292 17292 16348
rect 17228 16288 17292 16292
rect 17308 16348 17372 16352
rect 17308 16292 17312 16348
rect 17312 16292 17368 16348
rect 17368 16292 17372 16348
rect 17308 16288 17372 16292
rect 17388 16348 17452 16352
rect 17388 16292 17392 16348
rect 17392 16292 17448 16348
rect 17448 16292 17452 16348
rect 17388 16288 17452 16292
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 3831 15260 3895 15264
rect 3831 15204 3835 15260
rect 3835 15204 3891 15260
rect 3891 15204 3895 15260
rect 3831 15200 3895 15204
rect 3911 15260 3975 15264
rect 3911 15204 3915 15260
rect 3915 15204 3971 15260
rect 3971 15204 3975 15260
rect 3911 15200 3975 15204
rect 3991 15260 4055 15264
rect 3991 15204 3995 15260
rect 3995 15204 4051 15260
rect 4051 15204 4055 15260
rect 3991 15200 4055 15204
rect 4071 15260 4135 15264
rect 4071 15204 4075 15260
rect 4075 15204 4131 15260
rect 4131 15204 4135 15260
rect 4071 15200 4135 15204
rect 8270 15260 8334 15264
rect 8270 15204 8274 15260
rect 8274 15204 8330 15260
rect 8330 15204 8334 15260
rect 8270 15200 8334 15204
rect 8350 15260 8414 15264
rect 8350 15204 8354 15260
rect 8354 15204 8410 15260
rect 8410 15204 8414 15260
rect 8350 15200 8414 15204
rect 8430 15260 8494 15264
rect 8430 15204 8434 15260
rect 8434 15204 8490 15260
rect 8490 15204 8494 15260
rect 8430 15200 8494 15204
rect 8510 15260 8574 15264
rect 8510 15204 8514 15260
rect 8514 15204 8570 15260
rect 8570 15204 8574 15260
rect 8510 15200 8574 15204
rect 12709 15260 12773 15264
rect 12709 15204 12713 15260
rect 12713 15204 12769 15260
rect 12769 15204 12773 15260
rect 12709 15200 12773 15204
rect 12789 15260 12853 15264
rect 12789 15204 12793 15260
rect 12793 15204 12849 15260
rect 12849 15204 12853 15260
rect 12789 15200 12853 15204
rect 12869 15260 12933 15264
rect 12869 15204 12873 15260
rect 12873 15204 12929 15260
rect 12929 15204 12933 15260
rect 12869 15200 12933 15204
rect 12949 15260 13013 15264
rect 12949 15204 12953 15260
rect 12953 15204 13009 15260
rect 13009 15204 13013 15260
rect 12949 15200 13013 15204
rect 17148 15260 17212 15264
rect 17148 15204 17152 15260
rect 17152 15204 17208 15260
rect 17208 15204 17212 15260
rect 17148 15200 17212 15204
rect 17228 15260 17292 15264
rect 17228 15204 17232 15260
rect 17232 15204 17288 15260
rect 17288 15204 17292 15260
rect 17228 15200 17292 15204
rect 17308 15260 17372 15264
rect 17308 15204 17312 15260
rect 17312 15204 17368 15260
rect 17368 15204 17372 15260
rect 17308 15200 17372 15204
rect 17388 15260 17452 15264
rect 17388 15204 17392 15260
rect 17392 15204 17448 15260
rect 17448 15204 17452 15260
rect 17388 15200 17452 15204
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 3831 14172 3895 14176
rect 3831 14116 3835 14172
rect 3835 14116 3891 14172
rect 3891 14116 3895 14172
rect 3831 14112 3895 14116
rect 3911 14172 3975 14176
rect 3911 14116 3915 14172
rect 3915 14116 3971 14172
rect 3971 14116 3975 14172
rect 3911 14112 3975 14116
rect 3991 14172 4055 14176
rect 3991 14116 3995 14172
rect 3995 14116 4051 14172
rect 4051 14116 4055 14172
rect 3991 14112 4055 14116
rect 4071 14172 4135 14176
rect 4071 14116 4075 14172
rect 4075 14116 4131 14172
rect 4131 14116 4135 14172
rect 4071 14112 4135 14116
rect 8270 14172 8334 14176
rect 8270 14116 8274 14172
rect 8274 14116 8330 14172
rect 8330 14116 8334 14172
rect 8270 14112 8334 14116
rect 8350 14172 8414 14176
rect 8350 14116 8354 14172
rect 8354 14116 8410 14172
rect 8410 14116 8414 14172
rect 8350 14112 8414 14116
rect 8430 14172 8494 14176
rect 8430 14116 8434 14172
rect 8434 14116 8490 14172
rect 8490 14116 8494 14172
rect 8430 14112 8494 14116
rect 8510 14172 8574 14176
rect 8510 14116 8514 14172
rect 8514 14116 8570 14172
rect 8570 14116 8574 14172
rect 8510 14112 8574 14116
rect 12709 14172 12773 14176
rect 12709 14116 12713 14172
rect 12713 14116 12769 14172
rect 12769 14116 12773 14172
rect 12709 14112 12773 14116
rect 12789 14172 12853 14176
rect 12789 14116 12793 14172
rect 12793 14116 12849 14172
rect 12849 14116 12853 14172
rect 12789 14112 12853 14116
rect 12869 14172 12933 14176
rect 12869 14116 12873 14172
rect 12873 14116 12929 14172
rect 12929 14116 12933 14172
rect 12869 14112 12933 14116
rect 12949 14172 13013 14176
rect 12949 14116 12953 14172
rect 12953 14116 13009 14172
rect 13009 14116 13013 14172
rect 12949 14112 13013 14116
rect 17148 14172 17212 14176
rect 17148 14116 17152 14172
rect 17152 14116 17208 14172
rect 17208 14116 17212 14172
rect 17148 14112 17212 14116
rect 17228 14172 17292 14176
rect 17228 14116 17232 14172
rect 17232 14116 17288 14172
rect 17288 14116 17292 14172
rect 17228 14112 17292 14116
rect 17308 14172 17372 14176
rect 17308 14116 17312 14172
rect 17312 14116 17368 14172
rect 17368 14116 17372 14172
rect 17308 14112 17372 14116
rect 17388 14172 17452 14176
rect 17388 14116 17392 14172
rect 17392 14116 17448 14172
rect 17448 14116 17452 14172
rect 17388 14112 17452 14116
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 3831 13084 3895 13088
rect 3831 13028 3835 13084
rect 3835 13028 3891 13084
rect 3891 13028 3895 13084
rect 3831 13024 3895 13028
rect 3911 13084 3975 13088
rect 3911 13028 3915 13084
rect 3915 13028 3971 13084
rect 3971 13028 3975 13084
rect 3911 13024 3975 13028
rect 3991 13084 4055 13088
rect 3991 13028 3995 13084
rect 3995 13028 4051 13084
rect 4051 13028 4055 13084
rect 3991 13024 4055 13028
rect 4071 13084 4135 13088
rect 4071 13028 4075 13084
rect 4075 13028 4131 13084
rect 4131 13028 4135 13084
rect 4071 13024 4135 13028
rect 8270 13084 8334 13088
rect 8270 13028 8274 13084
rect 8274 13028 8330 13084
rect 8330 13028 8334 13084
rect 8270 13024 8334 13028
rect 8350 13084 8414 13088
rect 8350 13028 8354 13084
rect 8354 13028 8410 13084
rect 8410 13028 8414 13084
rect 8350 13024 8414 13028
rect 8430 13084 8494 13088
rect 8430 13028 8434 13084
rect 8434 13028 8490 13084
rect 8490 13028 8494 13084
rect 8430 13024 8494 13028
rect 8510 13084 8574 13088
rect 8510 13028 8514 13084
rect 8514 13028 8570 13084
rect 8570 13028 8574 13084
rect 8510 13024 8574 13028
rect 12709 13084 12773 13088
rect 12709 13028 12713 13084
rect 12713 13028 12769 13084
rect 12769 13028 12773 13084
rect 12709 13024 12773 13028
rect 12789 13084 12853 13088
rect 12789 13028 12793 13084
rect 12793 13028 12849 13084
rect 12849 13028 12853 13084
rect 12789 13024 12853 13028
rect 12869 13084 12933 13088
rect 12869 13028 12873 13084
rect 12873 13028 12929 13084
rect 12929 13028 12933 13084
rect 12869 13024 12933 13028
rect 12949 13084 13013 13088
rect 12949 13028 12953 13084
rect 12953 13028 13009 13084
rect 13009 13028 13013 13084
rect 12949 13024 13013 13028
rect 17148 13084 17212 13088
rect 17148 13028 17152 13084
rect 17152 13028 17208 13084
rect 17208 13028 17212 13084
rect 17148 13024 17212 13028
rect 17228 13084 17292 13088
rect 17228 13028 17232 13084
rect 17232 13028 17288 13084
rect 17288 13028 17292 13084
rect 17228 13024 17292 13028
rect 17308 13084 17372 13088
rect 17308 13028 17312 13084
rect 17312 13028 17368 13084
rect 17368 13028 17372 13084
rect 17308 13024 17372 13028
rect 17388 13084 17452 13088
rect 17388 13028 17392 13084
rect 17392 13028 17448 13084
rect 17448 13028 17452 13084
rect 17388 13024 17452 13028
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 3831 11996 3895 12000
rect 3831 11940 3835 11996
rect 3835 11940 3891 11996
rect 3891 11940 3895 11996
rect 3831 11936 3895 11940
rect 3911 11996 3975 12000
rect 3911 11940 3915 11996
rect 3915 11940 3971 11996
rect 3971 11940 3975 11996
rect 3911 11936 3975 11940
rect 3991 11996 4055 12000
rect 3991 11940 3995 11996
rect 3995 11940 4051 11996
rect 4051 11940 4055 11996
rect 3991 11936 4055 11940
rect 4071 11996 4135 12000
rect 4071 11940 4075 11996
rect 4075 11940 4131 11996
rect 4131 11940 4135 11996
rect 4071 11936 4135 11940
rect 8270 11996 8334 12000
rect 8270 11940 8274 11996
rect 8274 11940 8330 11996
rect 8330 11940 8334 11996
rect 8270 11936 8334 11940
rect 8350 11996 8414 12000
rect 8350 11940 8354 11996
rect 8354 11940 8410 11996
rect 8410 11940 8414 11996
rect 8350 11936 8414 11940
rect 8430 11996 8494 12000
rect 8430 11940 8434 11996
rect 8434 11940 8490 11996
rect 8490 11940 8494 11996
rect 8430 11936 8494 11940
rect 8510 11996 8574 12000
rect 8510 11940 8514 11996
rect 8514 11940 8570 11996
rect 8570 11940 8574 11996
rect 8510 11936 8574 11940
rect 12709 11996 12773 12000
rect 12709 11940 12713 11996
rect 12713 11940 12769 11996
rect 12769 11940 12773 11996
rect 12709 11936 12773 11940
rect 12789 11996 12853 12000
rect 12789 11940 12793 11996
rect 12793 11940 12849 11996
rect 12849 11940 12853 11996
rect 12789 11936 12853 11940
rect 12869 11996 12933 12000
rect 12869 11940 12873 11996
rect 12873 11940 12929 11996
rect 12929 11940 12933 11996
rect 12869 11936 12933 11940
rect 12949 11996 13013 12000
rect 12949 11940 12953 11996
rect 12953 11940 13009 11996
rect 13009 11940 13013 11996
rect 12949 11936 13013 11940
rect 17148 11996 17212 12000
rect 17148 11940 17152 11996
rect 17152 11940 17208 11996
rect 17208 11940 17212 11996
rect 17148 11936 17212 11940
rect 17228 11996 17292 12000
rect 17228 11940 17232 11996
rect 17232 11940 17288 11996
rect 17288 11940 17292 11996
rect 17228 11936 17292 11940
rect 17308 11996 17372 12000
rect 17308 11940 17312 11996
rect 17312 11940 17368 11996
rect 17368 11940 17372 11996
rect 17308 11936 17372 11940
rect 17388 11996 17452 12000
rect 17388 11940 17392 11996
rect 17392 11940 17448 11996
rect 17448 11940 17452 11996
rect 17388 11936 17452 11940
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 3831 10908 3895 10912
rect 3831 10852 3835 10908
rect 3835 10852 3891 10908
rect 3891 10852 3895 10908
rect 3831 10848 3895 10852
rect 3911 10908 3975 10912
rect 3911 10852 3915 10908
rect 3915 10852 3971 10908
rect 3971 10852 3975 10908
rect 3911 10848 3975 10852
rect 3991 10908 4055 10912
rect 3991 10852 3995 10908
rect 3995 10852 4051 10908
rect 4051 10852 4055 10908
rect 3991 10848 4055 10852
rect 4071 10908 4135 10912
rect 4071 10852 4075 10908
rect 4075 10852 4131 10908
rect 4131 10852 4135 10908
rect 4071 10848 4135 10852
rect 8270 10908 8334 10912
rect 8270 10852 8274 10908
rect 8274 10852 8330 10908
rect 8330 10852 8334 10908
rect 8270 10848 8334 10852
rect 8350 10908 8414 10912
rect 8350 10852 8354 10908
rect 8354 10852 8410 10908
rect 8410 10852 8414 10908
rect 8350 10848 8414 10852
rect 8430 10908 8494 10912
rect 8430 10852 8434 10908
rect 8434 10852 8490 10908
rect 8490 10852 8494 10908
rect 8430 10848 8494 10852
rect 8510 10908 8574 10912
rect 8510 10852 8514 10908
rect 8514 10852 8570 10908
rect 8570 10852 8574 10908
rect 8510 10848 8574 10852
rect 12709 10908 12773 10912
rect 12709 10852 12713 10908
rect 12713 10852 12769 10908
rect 12769 10852 12773 10908
rect 12709 10848 12773 10852
rect 12789 10908 12853 10912
rect 12789 10852 12793 10908
rect 12793 10852 12849 10908
rect 12849 10852 12853 10908
rect 12789 10848 12853 10852
rect 12869 10908 12933 10912
rect 12869 10852 12873 10908
rect 12873 10852 12929 10908
rect 12929 10852 12933 10908
rect 12869 10848 12933 10852
rect 12949 10908 13013 10912
rect 12949 10852 12953 10908
rect 12953 10852 13009 10908
rect 13009 10852 13013 10908
rect 12949 10848 13013 10852
rect 17148 10908 17212 10912
rect 17148 10852 17152 10908
rect 17152 10852 17208 10908
rect 17208 10852 17212 10908
rect 17148 10848 17212 10852
rect 17228 10908 17292 10912
rect 17228 10852 17232 10908
rect 17232 10852 17288 10908
rect 17288 10852 17292 10908
rect 17228 10848 17292 10852
rect 17308 10908 17372 10912
rect 17308 10852 17312 10908
rect 17312 10852 17368 10908
rect 17368 10852 17372 10908
rect 17308 10848 17372 10852
rect 17388 10908 17452 10912
rect 17388 10852 17392 10908
rect 17392 10852 17448 10908
rect 17448 10852 17452 10908
rect 17388 10848 17452 10852
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 3831 9820 3895 9824
rect 3831 9764 3835 9820
rect 3835 9764 3891 9820
rect 3891 9764 3895 9820
rect 3831 9760 3895 9764
rect 3911 9820 3975 9824
rect 3911 9764 3915 9820
rect 3915 9764 3971 9820
rect 3971 9764 3975 9820
rect 3911 9760 3975 9764
rect 3991 9820 4055 9824
rect 3991 9764 3995 9820
rect 3995 9764 4051 9820
rect 4051 9764 4055 9820
rect 3991 9760 4055 9764
rect 4071 9820 4135 9824
rect 4071 9764 4075 9820
rect 4075 9764 4131 9820
rect 4131 9764 4135 9820
rect 4071 9760 4135 9764
rect 8270 9820 8334 9824
rect 8270 9764 8274 9820
rect 8274 9764 8330 9820
rect 8330 9764 8334 9820
rect 8270 9760 8334 9764
rect 8350 9820 8414 9824
rect 8350 9764 8354 9820
rect 8354 9764 8410 9820
rect 8410 9764 8414 9820
rect 8350 9760 8414 9764
rect 8430 9820 8494 9824
rect 8430 9764 8434 9820
rect 8434 9764 8490 9820
rect 8490 9764 8494 9820
rect 8430 9760 8494 9764
rect 8510 9820 8574 9824
rect 8510 9764 8514 9820
rect 8514 9764 8570 9820
rect 8570 9764 8574 9820
rect 8510 9760 8574 9764
rect 12709 9820 12773 9824
rect 12709 9764 12713 9820
rect 12713 9764 12769 9820
rect 12769 9764 12773 9820
rect 12709 9760 12773 9764
rect 12789 9820 12853 9824
rect 12789 9764 12793 9820
rect 12793 9764 12849 9820
rect 12849 9764 12853 9820
rect 12789 9760 12853 9764
rect 12869 9820 12933 9824
rect 12869 9764 12873 9820
rect 12873 9764 12929 9820
rect 12929 9764 12933 9820
rect 12869 9760 12933 9764
rect 12949 9820 13013 9824
rect 12949 9764 12953 9820
rect 12953 9764 13009 9820
rect 13009 9764 13013 9820
rect 12949 9760 13013 9764
rect 17148 9820 17212 9824
rect 17148 9764 17152 9820
rect 17152 9764 17208 9820
rect 17208 9764 17212 9820
rect 17148 9760 17212 9764
rect 17228 9820 17292 9824
rect 17228 9764 17232 9820
rect 17232 9764 17288 9820
rect 17288 9764 17292 9820
rect 17228 9760 17292 9764
rect 17308 9820 17372 9824
rect 17308 9764 17312 9820
rect 17312 9764 17368 9820
rect 17368 9764 17372 9820
rect 17308 9760 17372 9764
rect 17388 9820 17452 9824
rect 17388 9764 17392 9820
rect 17392 9764 17448 9820
rect 17448 9764 17452 9820
rect 17388 9760 17452 9764
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 3831 8732 3895 8736
rect 3831 8676 3835 8732
rect 3835 8676 3891 8732
rect 3891 8676 3895 8732
rect 3831 8672 3895 8676
rect 3911 8732 3975 8736
rect 3911 8676 3915 8732
rect 3915 8676 3971 8732
rect 3971 8676 3975 8732
rect 3911 8672 3975 8676
rect 3991 8732 4055 8736
rect 3991 8676 3995 8732
rect 3995 8676 4051 8732
rect 4051 8676 4055 8732
rect 3991 8672 4055 8676
rect 4071 8732 4135 8736
rect 4071 8676 4075 8732
rect 4075 8676 4131 8732
rect 4131 8676 4135 8732
rect 4071 8672 4135 8676
rect 8270 8732 8334 8736
rect 8270 8676 8274 8732
rect 8274 8676 8330 8732
rect 8330 8676 8334 8732
rect 8270 8672 8334 8676
rect 8350 8732 8414 8736
rect 8350 8676 8354 8732
rect 8354 8676 8410 8732
rect 8410 8676 8414 8732
rect 8350 8672 8414 8676
rect 8430 8732 8494 8736
rect 8430 8676 8434 8732
rect 8434 8676 8490 8732
rect 8490 8676 8494 8732
rect 8430 8672 8494 8676
rect 8510 8732 8574 8736
rect 8510 8676 8514 8732
rect 8514 8676 8570 8732
rect 8570 8676 8574 8732
rect 8510 8672 8574 8676
rect 12709 8732 12773 8736
rect 12709 8676 12713 8732
rect 12713 8676 12769 8732
rect 12769 8676 12773 8732
rect 12709 8672 12773 8676
rect 12789 8732 12853 8736
rect 12789 8676 12793 8732
rect 12793 8676 12849 8732
rect 12849 8676 12853 8732
rect 12789 8672 12853 8676
rect 12869 8732 12933 8736
rect 12869 8676 12873 8732
rect 12873 8676 12929 8732
rect 12929 8676 12933 8732
rect 12869 8672 12933 8676
rect 12949 8732 13013 8736
rect 12949 8676 12953 8732
rect 12953 8676 13009 8732
rect 13009 8676 13013 8732
rect 12949 8672 13013 8676
rect 17148 8732 17212 8736
rect 17148 8676 17152 8732
rect 17152 8676 17208 8732
rect 17208 8676 17212 8732
rect 17148 8672 17212 8676
rect 17228 8732 17292 8736
rect 17228 8676 17232 8732
rect 17232 8676 17288 8732
rect 17288 8676 17292 8732
rect 17228 8672 17292 8676
rect 17308 8732 17372 8736
rect 17308 8676 17312 8732
rect 17312 8676 17368 8732
rect 17368 8676 17372 8732
rect 17308 8672 17372 8676
rect 17388 8732 17452 8736
rect 17388 8676 17392 8732
rect 17392 8676 17448 8732
rect 17448 8676 17452 8732
rect 17388 8672 17452 8676
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 3831 7644 3895 7648
rect 3831 7588 3835 7644
rect 3835 7588 3891 7644
rect 3891 7588 3895 7644
rect 3831 7584 3895 7588
rect 3911 7644 3975 7648
rect 3911 7588 3915 7644
rect 3915 7588 3971 7644
rect 3971 7588 3975 7644
rect 3911 7584 3975 7588
rect 3991 7644 4055 7648
rect 3991 7588 3995 7644
rect 3995 7588 4051 7644
rect 4051 7588 4055 7644
rect 3991 7584 4055 7588
rect 4071 7644 4135 7648
rect 4071 7588 4075 7644
rect 4075 7588 4131 7644
rect 4131 7588 4135 7644
rect 4071 7584 4135 7588
rect 8270 7644 8334 7648
rect 8270 7588 8274 7644
rect 8274 7588 8330 7644
rect 8330 7588 8334 7644
rect 8270 7584 8334 7588
rect 8350 7644 8414 7648
rect 8350 7588 8354 7644
rect 8354 7588 8410 7644
rect 8410 7588 8414 7644
rect 8350 7584 8414 7588
rect 8430 7644 8494 7648
rect 8430 7588 8434 7644
rect 8434 7588 8490 7644
rect 8490 7588 8494 7644
rect 8430 7584 8494 7588
rect 8510 7644 8574 7648
rect 8510 7588 8514 7644
rect 8514 7588 8570 7644
rect 8570 7588 8574 7644
rect 8510 7584 8574 7588
rect 12709 7644 12773 7648
rect 12709 7588 12713 7644
rect 12713 7588 12769 7644
rect 12769 7588 12773 7644
rect 12709 7584 12773 7588
rect 12789 7644 12853 7648
rect 12789 7588 12793 7644
rect 12793 7588 12849 7644
rect 12849 7588 12853 7644
rect 12789 7584 12853 7588
rect 12869 7644 12933 7648
rect 12869 7588 12873 7644
rect 12873 7588 12929 7644
rect 12929 7588 12933 7644
rect 12869 7584 12933 7588
rect 12949 7644 13013 7648
rect 12949 7588 12953 7644
rect 12953 7588 13009 7644
rect 13009 7588 13013 7644
rect 12949 7584 13013 7588
rect 17148 7644 17212 7648
rect 17148 7588 17152 7644
rect 17152 7588 17208 7644
rect 17208 7588 17212 7644
rect 17148 7584 17212 7588
rect 17228 7644 17292 7648
rect 17228 7588 17232 7644
rect 17232 7588 17288 7644
rect 17288 7588 17292 7644
rect 17228 7584 17292 7588
rect 17308 7644 17372 7648
rect 17308 7588 17312 7644
rect 17312 7588 17368 7644
rect 17368 7588 17372 7644
rect 17308 7584 17372 7588
rect 17388 7644 17452 7648
rect 17388 7588 17392 7644
rect 17392 7588 17448 7644
rect 17448 7588 17452 7644
rect 17388 7584 17452 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 3831 6556 3895 6560
rect 3831 6500 3835 6556
rect 3835 6500 3891 6556
rect 3891 6500 3895 6556
rect 3831 6496 3895 6500
rect 3911 6556 3975 6560
rect 3911 6500 3915 6556
rect 3915 6500 3971 6556
rect 3971 6500 3975 6556
rect 3911 6496 3975 6500
rect 3991 6556 4055 6560
rect 3991 6500 3995 6556
rect 3995 6500 4051 6556
rect 4051 6500 4055 6556
rect 3991 6496 4055 6500
rect 4071 6556 4135 6560
rect 4071 6500 4075 6556
rect 4075 6500 4131 6556
rect 4131 6500 4135 6556
rect 4071 6496 4135 6500
rect 8270 6556 8334 6560
rect 8270 6500 8274 6556
rect 8274 6500 8330 6556
rect 8330 6500 8334 6556
rect 8270 6496 8334 6500
rect 8350 6556 8414 6560
rect 8350 6500 8354 6556
rect 8354 6500 8410 6556
rect 8410 6500 8414 6556
rect 8350 6496 8414 6500
rect 8430 6556 8494 6560
rect 8430 6500 8434 6556
rect 8434 6500 8490 6556
rect 8490 6500 8494 6556
rect 8430 6496 8494 6500
rect 8510 6556 8574 6560
rect 8510 6500 8514 6556
rect 8514 6500 8570 6556
rect 8570 6500 8574 6556
rect 8510 6496 8574 6500
rect 12709 6556 12773 6560
rect 12709 6500 12713 6556
rect 12713 6500 12769 6556
rect 12769 6500 12773 6556
rect 12709 6496 12773 6500
rect 12789 6556 12853 6560
rect 12789 6500 12793 6556
rect 12793 6500 12849 6556
rect 12849 6500 12853 6556
rect 12789 6496 12853 6500
rect 12869 6556 12933 6560
rect 12869 6500 12873 6556
rect 12873 6500 12929 6556
rect 12929 6500 12933 6556
rect 12869 6496 12933 6500
rect 12949 6556 13013 6560
rect 12949 6500 12953 6556
rect 12953 6500 13009 6556
rect 13009 6500 13013 6556
rect 12949 6496 13013 6500
rect 17148 6556 17212 6560
rect 17148 6500 17152 6556
rect 17152 6500 17208 6556
rect 17208 6500 17212 6556
rect 17148 6496 17212 6500
rect 17228 6556 17292 6560
rect 17228 6500 17232 6556
rect 17232 6500 17288 6556
rect 17288 6500 17292 6556
rect 17228 6496 17292 6500
rect 17308 6556 17372 6560
rect 17308 6500 17312 6556
rect 17312 6500 17368 6556
rect 17368 6500 17372 6556
rect 17308 6496 17372 6500
rect 17388 6556 17452 6560
rect 17388 6500 17392 6556
rect 17392 6500 17448 6556
rect 17448 6500 17452 6556
rect 17388 6496 17452 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 3831 5468 3895 5472
rect 3831 5412 3835 5468
rect 3835 5412 3891 5468
rect 3891 5412 3895 5468
rect 3831 5408 3895 5412
rect 3911 5468 3975 5472
rect 3911 5412 3915 5468
rect 3915 5412 3971 5468
rect 3971 5412 3975 5468
rect 3911 5408 3975 5412
rect 3991 5468 4055 5472
rect 3991 5412 3995 5468
rect 3995 5412 4051 5468
rect 4051 5412 4055 5468
rect 3991 5408 4055 5412
rect 4071 5468 4135 5472
rect 4071 5412 4075 5468
rect 4075 5412 4131 5468
rect 4131 5412 4135 5468
rect 4071 5408 4135 5412
rect 8270 5468 8334 5472
rect 8270 5412 8274 5468
rect 8274 5412 8330 5468
rect 8330 5412 8334 5468
rect 8270 5408 8334 5412
rect 8350 5468 8414 5472
rect 8350 5412 8354 5468
rect 8354 5412 8410 5468
rect 8410 5412 8414 5468
rect 8350 5408 8414 5412
rect 8430 5468 8494 5472
rect 8430 5412 8434 5468
rect 8434 5412 8490 5468
rect 8490 5412 8494 5468
rect 8430 5408 8494 5412
rect 8510 5468 8574 5472
rect 8510 5412 8514 5468
rect 8514 5412 8570 5468
rect 8570 5412 8574 5468
rect 8510 5408 8574 5412
rect 12709 5468 12773 5472
rect 12709 5412 12713 5468
rect 12713 5412 12769 5468
rect 12769 5412 12773 5468
rect 12709 5408 12773 5412
rect 12789 5468 12853 5472
rect 12789 5412 12793 5468
rect 12793 5412 12849 5468
rect 12849 5412 12853 5468
rect 12789 5408 12853 5412
rect 12869 5468 12933 5472
rect 12869 5412 12873 5468
rect 12873 5412 12929 5468
rect 12929 5412 12933 5468
rect 12869 5408 12933 5412
rect 12949 5468 13013 5472
rect 12949 5412 12953 5468
rect 12953 5412 13009 5468
rect 13009 5412 13013 5468
rect 12949 5408 13013 5412
rect 17148 5468 17212 5472
rect 17148 5412 17152 5468
rect 17152 5412 17208 5468
rect 17208 5412 17212 5468
rect 17148 5408 17212 5412
rect 17228 5468 17292 5472
rect 17228 5412 17232 5468
rect 17232 5412 17288 5468
rect 17288 5412 17292 5468
rect 17228 5408 17292 5412
rect 17308 5468 17372 5472
rect 17308 5412 17312 5468
rect 17312 5412 17368 5468
rect 17368 5412 17372 5468
rect 17308 5408 17372 5412
rect 17388 5468 17452 5472
rect 17388 5412 17392 5468
rect 17392 5412 17448 5468
rect 17448 5412 17452 5468
rect 17388 5408 17452 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 3831 4380 3895 4384
rect 3831 4324 3835 4380
rect 3835 4324 3891 4380
rect 3891 4324 3895 4380
rect 3831 4320 3895 4324
rect 3911 4380 3975 4384
rect 3911 4324 3915 4380
rect 3915 4324 3971 4380
rect 3971 4324 3975 4380
rect 3911 4320 3975 4324
rect 3991 4380 4055 4384
rect 3991 4324 3995 4380
rect 3995 4324 4051 4380
rect 4051 4324 4055 4380
rect 3991 4320 4055 4324
rect 4071 4380 4135 4384
rect 4071 4324 4075 4380
rect 4075 4324 4131 4380
rect 4131 4324 4135 4380
rect 4071 4320 4135 4324
rect 8270 4380 8334 4384
rect 8270 4324 8274 4380
rect 8274 4324 8330 4380
rect 8330 4324 8334 4380
rect 8270 4320 8334 4324
rect 8350 4380 8414 4384
rect 8350 4324 8354 4380
rect 8354 4324 8410 4380
rect 8410 4324 8414 4380
rect 8350 4320 8414 4324
rect 8430 4380 8494 4384
rect 8430 4324 8434 4380
rect 8434 4324 8490 4380
rect 8490 4324 8494 4380
rect 8430 4320 8494 4324
rect 8510 4380 8574 4384
rect 8510 4324 8514 4380
rect 8514 4324 8570 4380
rect 8570 4324 8574 4380
rect 8510 4320 8574 4324
rect 12709 4380 12773 4384
rect 12709 4324 12713 4380
rect 12713 4324 12769 4380
rect 12769 4324 12773 4380
rect 12709 4320 12773 4324
rect 12789 4380 12853 4384
rect 12789 4324 12793 4380
rect 12793 4324 12849 4380
rect 12849 4324 12853 4380
rect 12789 4320 12853 4324
rect 12869 4380 12933 4384
rect 12869 4324 12873 4380
rect 12873 4324 12929 4380
rect 12929 4324 12933 4380
rect 12869 4320 12933 4324
rect 12949 4380 13013 4384
rect 12949 4324 12953 4380
rect 12953 4324 13009 4380
rect 13009 4324 13013 4380
rect 12949 4320 13013 4324
rect 17148 4380 17212 4384
rect 17148 4324 17152 4380
rect 17152 4324 17208 4380
rect 17208 4324 17212 4380
rect 17148 4320 17212 4324
rect 17228 4380 17292 4384
rect 17228 4324 17232 4380
rect 17232 4324 17288 4380
rect 17288 4324 17292 4380
rect 17228 4320 17292 4324
rect 17308 4380 17372 4384
rect 17308 4324 17312 4380
rect 17312 4324 17368 4380
rect 17368 4324 17372 4380
rect 17308 4320 17372 4324
rect 17388 4380 17452 4384
rect 17388 4324 17392 4380
rect 17392 4324 17448 4380
rect 17448 4324 17452 4380
rect 17388 4320 17452 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 3831 3292 3895 3296
rect 3831 3236 3835 3292
rect 3835 3236 3891 3292
rect 3891 3236 3895 3292
rect 3831 3232 3895 3236
rect 3911 3292 3975 3296
rect 3911 3236 3915 3292
rect 3915 3236 3971 3292
rect 3971 3236 3975 3292
rect 3911 3232 3975 3236
rect 3991 3292 4055 3296
rect 3991 3236 3995 3292
rect 3995 3236 4051 3292
rect 4051 3236 4055 3292
rect 3991 3232 4055 3236
rect 4071 3292 4135 3296
rect 4071 3236 4075 3292
rect 4075 3236 4131 3292
rect 4131 3236 4135 3292
rect 4071 3232 4135 3236
rect 8270 3292 8334 3296
rect 8270 3236 8274 3292
rect 8274 3236 8330 3292
rect 8330 3236 8334 3292
rect 8270 3232 8334 3236
rect 8350 3292 8414 3296
rect 8350 3236 8354 3292
rect 8354 3236 8410 3292
rect 8410 3236 8414 3292
rect 8350 3232 8414 3236
rect 8430 3292 8494 3296
rect 8430 3236 8434 3292
rect 8434 3236 8490 3292
rect 8490 3236 8494 3292
rect 8430 3232 8494 3236
rect 8510 3292 8574 3296
rect 8510 3236 8514 3292
rect 8514 3236 8570 3292
rect 8570 3236 8574 3292
rect 8510 3232 8574 3236
rect 12709 3292 12773 3296
rect 12709 3236 12713 3292
rect 12713 3236 12769 3292
rect 12769 3236 12773 3292
rect 12709 3232 12773 3236
rect 12789 3292 12853 3296
rect 12789 3236 12793 3292
rect 12793 3236 12849 3292
rect 12849 3236 12853 3292
rect 12789 3232 12853 3236
rect 12869 3292 12933 3296
rect 12869 3236 12873 3292
rect 12873 3236 12929 3292
rect 12929 3236 12933 3292
rect 12869 3232 12933 3236
rect 12949 3292 13013 3296
rect 12949 3236 12953 3292
rect 12953 3236 13009 3292
rect 13009 3236 13013 3292
rect 12949 3232 13013 3236
rect 17148 3292 17212 3296
rect 17148 3236 17152 3292
rect 17152 3236 17208 3292
rect 17208 3236 17212 3292
rect 17148 3232 17212 3236
rect 17228 3292 17292 3296
rect 17228 3236 17232 3292
rect 17232 3236 17288 3292
rect 17288 3236 17292 3292
rect 17228 3232 17292 3236
rect 17308 3292 17372 3296
rect 17308 3236 17312 3292
rect 17312 3236 17368 3292
rect 17368 3236 17372 3292
rect 17308 3232 17372 3236
rect 17388 3292 17452 3296
rect 17388 3236 17392 3292
rect 17392 3236 17448 3292
rect 17448 3236 17452 3292
rect 17388 3232 17452 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 3831 2204 3895 2208
rect 3831 2148 3835 2204
rect 3835 2148 3891 2204
rect 3891 2148 3895 2204
rect 3831 2144 3895 2148
rect 3911 2204 3975 2208
rect 3911 2148 3915 2204
rect 3915 2148 3971 2204
rect 3971 2148 3975 2204
rect 3911 2144 3975 2148
rect 3991 2204 4055 2208
rect 3991 2148 3995 2204
rect 3995 2148 4051 2204
rect 4051 2148 4055 2204
rect 3991 2144 4055 2148
rect 4071 2204 4135 2208
rect 4071 2148 4075 2204
rect 4075 2148 4131 2204
rect 4131 2148 4135 2204
rect 4071 2144 4135 2148
rect 8270 2204 8334 2208
rect 8270 2148 8274 2204
rect 8274 2148 8330 2204
rect 8330 2148 8334 2204
rect 8270 2144 8334 2148
rect 8350 2204 8414 2208
rect 8350 2148 8354 2204
rect 8354 2148 8410 2204
rect 8410 2148 8414 2204
rect 8350 2144 8414 2148
rect 8430 2204 8494 2208
rect 8430 2148 8434 2204
rect 8434 2148 8490 2204
rect 8490 2148 8494 2204
rect 8430 2144 8494 2148
rect 8510 2204 8574 2208
rect 8510 2148 8514 2204
rect 8514 2148 8570 2204
rect 8570 2148 8574 2204
rect 8510 2144 8574 2148
rect 12709 2204 12773 2208
rect 12709 2148 12713 2204
rect 12713 2148 12769 2204
rect 12769 2148 12773 2204
rect 12709 2144 12773 2148
rect 12789 2204 12853 2208
rect 12789 2148 12793 2204
rect 12793 2148 12849 2204
rect 12849 2148 12853 2204
rect 12789 2144 12853 2148
rect 12869 2204 12933 2208
rect 12869 2148 12873 2204
rect 12873 2148 12929 2204
rect 12929 2148 12933 2204
rect 12869 2144 12933 2148
rect 12949 2204 13013 2208
rect 12949 2148 12953 2204
rect 12953 2148 13009 2204
rect 13009 2148 13013 2204
rect 12949 2144 13013 2148
rect 17148 2204 17212 2208
rect 17148 2148 17152 2204
rect 17152 2148 17208 2204
rect 17208 2148 17212 2204
rect 17148 2144 17212 2148
rect 17228 2204 17292 2208
rect 17228 2148 17232 2204
rect 17232 2148 17288 2204
rect 17288 2148 17292 2204
rect 17228 2144 17292 2148
rect 17308 2204 17372 2208
rect 17308 2148 17312 2204
rect 17312 2148 17368 2204
rect 17368 2148 17372 2204
rect 17308 2144 17372 2148
rect 17388 2204 17452 2208
rect 17388 2148 17392 2204
rect 17392 2148 17448 2204
rect 17448 2148 17452 2204
rect 17388 2144 17452 2148
<< metal4 >>
rect 3163 16896 3483 17456
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3163 15808 3483 16832
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 15622 3483 15744
rect 3163 15386 3205 15622
rect 3441 15386 3483 15622
rect 3163 14720 3483 15386
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11814 3483 12480
rect 3163 11578 3205 11814
rect 3441 11578 3483 11814
rect 3163 11456 3483 11578
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 8006 3483 8128
rect 3163 7770 3205 8006
rect 3441 7770 3483 8006
rect 3163 7104 3483 7770
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 4198 3483 4864
rect 3163 3962 3205 4198
rect 3441 3962 3483 4198
rect 3163 3840 3483 3962
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 3823 17440 4143 17456
rect 3823 17376 3831 17440
rect 3895 17376 3911 17440
rect 3975 17376 3991 17440
rect 4055 17376 4071 17440
rect 4135 17376 4143 17440
rect 3823 16352 4143 17376
rect 3823 16288 3831 16352
rect 3895 16288 3911 16352
rect 3975 16288 3991 16352
rect 4055 16288 4071 16352
rect 4135 16288 4143 16352
rect 3823 16282 4143 16288
rect 3823 16046 3865 16282
rect 4101 16046 4143 16282
rect 3823 15264 4143 16046
rect 3823 15200 3831 15264
rect 3895 15200 3911 15264
rect 3975 15200 3991 15264
rect 4055 15200 4071 15264
rect 4135 15200 4143 15264
rect 3823 14176 4143 15200
rect 3823 14112 3831 14176
rect 3895 14112 3911 14176
rect 3975 14112 3991 14176
rect 4055 14112 4071 14176
rect 4135 14112 4143 14176
rect 3823 13088 4143 14112
rect 3823 13024 3831 13088
rect 3895 13024 3911 13088
rect 3975 13024 3991 13088
rect 4055 13024 4071 13088
rect 4135 13024 4143 13088
rect 3823 12474 4143 13024
rect 3823 12238 3865 12474
rect 4101 12238 4143 12474
rect 3823 12000 4143 12238
rect 3823 11936 3831 12000
rect 3895 11936 3911 12000
rect 3975 11936 3991 12000
rect 4055 11936 4071 12000
rect 4135 11936 4143 12000
rect 3823 10912 4143 11936
rect 3823 10848 3831 10912
rect 3895 10848 3911 10912
rect 3975 10848 3991 10912
rect 4055 10848 4071 10912
rect 4135 10848 4143 10912
rect 3823 9824 4143 10848
rect 3823 9760 3831 9824
rect 3895 9760 3911 9824
rect 3975 9760 3991 9824
rect 4055 9760 4071 9824
rect 4135 9760 4143 9824
rect 3823 8736 4143 9760
rect 3823 8672 3831 8736
rect 3895 8672 3911 8736
rect 3975 8672 3991 8736
rect 4055 8672 4071 8736
rect 4135 8672 4143 8736
rect 3823 8666 4143 8672
rect 3823 8430 3865 8666
rect 4101 8430 4143 8666
rect 3823 7648 4143 8430
rect 3823 7584 3831 7648
rect 3895 7584 3911 7648
rect 3975 7584 3991 7648
rect 4055 7584 4071 7648
rect 4135 7584 4143 7648
rect 3823 6560 4143 7584
rect 3823 6496 3831 6560
rect 3895 6496 3911 6560
rect 3975 6496 3991 6560
rect 4055 6496 4071 6560
rect 4135 6496 4143 6560
rect 3823 5472 4143 6496
rect 3823 5408 3831 5472
rect 3895 5408 3911 5472
rect 3975 5408 3991 5472
rect 4055 5408 4071 5472
rect 4135 5408 4143 5472
rect 3823 4858 4143 5408
rect 3823 4622 3865 4858
rect 4101 4622 4143 4858
rect 3823 4384 4143 4622
rect 3823 4320 3831 4384
rect 3895 4320 3911 4384
rect 3975 4320 3991 4384
rect 4055 4320 4071 4384
rect 4135 4320 4143 4384
rect 3823 3296 4143 4320
rect 3823 3232 3831 3296
rect 3895 3232 3911 3296
rect 3975 3232 3991 3296
rect 4055 3232 4071 3296
rect 4135 3232 4143 3296
rect 3823 2208 4143 3232
rect 3823 2144 3831 2208
rect 3895 2144 3911 2208
rect 3975 2144 3991 2208
rect 4055 2144 4071 2208
rect 4135 2144 4143 2208
rect 3823 2128 4143 2144
rect 7602 16896 7922 17456
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 15622 7922 15744
rect 7602 15386 7644 15622
rect 7880 15386 7922 15622
rect 7602 14720 7922 15386
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11814 7922 12480
rect 7602 11578 7644 11814
rect 7880 11578 7922 11814
rect 7602 11456 7922 11578
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 8006 7922 8128
rect 7602 7770 7644 8006
rect 7880 7770 7922 8006
rect 7602 7104 7922 7770
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 4198 7922 4864
rect 7602 3962 7644 4198
rect 7880 3962 7922 4198
rect 7602 3840 7922 3962
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 8262 17440 8582 17456
rect 8262 17376 8270 17440
rect 8334 17376 8350 17440
rect 8414 17376 8430 17440
rect 8494 17376 8510 17440
rect 8574 17376 8582 17440
rect 8262 16352 8582 17376
rect 8262 16288 8270 16352
rect 8334 16288 8350 16352
rect 8414 16288 8430 16352
rect 8494 16288 8510 16352
rect 8574 16288 8582 16352
rect 8262 16282 8582 16288
rect 8262 16046 8304 16282
rect 8540 16046 8582 16282
rect 8262 15264 8582 16046
rect 8262 15200 8270 15264
rect 8334 15200 8350 15264
rect 8414 15200 8430 15264
rect 8494 15200 8510 15264
rect 8574 15200 8582 15264
rect 8262 14176 8582 15200
rect 8262 14112 8270 14176
rect 8334 14112 8350 14176
rect 8414 14112 8430 14176
rect 8494 14112 8510 14176
rect 8574 14112 8582 14176
rect 8262 13088 8582 14112
rect 8262 13024 8270 13088
rect 8334 13024 8350 13088
rect 8414 13024 8430 13088
rect 8494 13024 8510 13088
rect 8574 13024 8582 13088
rect 8262 12474 8582 13024
rect 8262 12238 8304 12474
rect 8540 12238 8582 12474
rect 8262 12000 8582 12238
rect 8262 11936 8270 12000
rect 8334 11936 8350 12000
rect 8414 11936 8430 12000
rect 8494 11936 8510 12000
rect 8574 11936 8582 12000
rect 8262 10912 8582 11936
rect 8262 10848 8270 10912
rect 8334 10848 8350 10912
rect 8414 10848 8430 10912
rect 8494 10848 8510 10912
rect 8574 10848 8582 10912
rect 8262 9824 8582 10848
rect 8262 9760 8270 9824
rect 8334 9760 8350 9824
rect 8414 9760 8430 9824
rect 8494 9760 8510 9824
rect 8574 9760 8582 9824
rect 8262 8736 8582 9760
rect 8262 8672 8270 8736
rect 8334 8672 8350 8736
rect 8414 8672 8430 8736
rect 8494 8672 8510 8736
rect 8574 8672 8582 8736
rect 8262 8666 8582 8672
rect 8262 8430 8304 8666
rect 8540 8430 8582 8666
rect 8262 7648 8582 8430
rect 8262 7584 8270 7648
rect 8334 7584 8350 7648
rect 8414 7584 8430 7648
rect 8494 7584 8510 7648
rect 8574 7584 8582 7648
rect 8262 6560 8582 7584
rect 8262 6496 8270 6560
rect 8334 6496 8350 6560
rect 8414 6496 8430 6560
rect 8494 6496 8510 6560
rect 8574 6496 8582 6560
rect 8262 5472 8582 6496
rect 8262 5408 8270 5472
rect 8334 5408 8350 5472
rect 8414 5408 8430 5472
rect 8494 5408 8510 5472
rect 8574 5408 8582 5472
rect 8262 4858 8582 5408
rect 8262 4622 8304 4858
rect 8540 4622 8582 4858
rect 8262 4384 8582 4622
rect 8262 4320 8270 4384
rect 8334 4320 8350 4384
rect 8414 4320 8430 4384
rect 8494 4320 8510 4384
rect 8574 4320 8582 4384
rect 8262 3296 8582 4320
rect 8262 3232 8270 3296
rect 8334 3232 8350 3296
rect 8414 3232 8430 3296
rect 8494 3232 8510 3296
rect 8574 3232 8582 3296
rect 8262 2208 8582 3232
rect 8262 2144 8270 2208
rect 8334 2144 8350 2208
rect 8414 2144 8430 2208
rect 8494 2144 8510 2208
rect 8574 2144 8582 2208
rect 8262 2128 8582 2144
rect 12041 16896 12361 17456
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 15622 12361 15744
rect 12041 15386 12083 15622
rect 12319 15386 12361 15622
rect 12041 14720 12361 15386
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11814 12361 12480
rect 12041 11578 12083 11814
rect 12319 11578 12361 11814
rect 12041 11456 12361 11578
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 8006 12361 8128
rect 12041 7770 12083 8006
rect 12319 7770 12361 8006
rect 12041 7104 12361 7770
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 4198 12361 4864
rect 12041 3962 12083 4198
rect 12319 3962 12361 4198
rect 12041 3840 12361 3962
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 12701 17440 13021 17456
rect 12701 17376 12709 17440
rect 12773 17376 12789 17440
rect 12853 17376 12869 17440
rect 12933 17376 12949 17440
rect 13013 17376 13021 17440
rect 12701 16352 13021 17376
rect 12701 16288 12709 16352
rect 12773 16288 12789 16352
rect 12853 16288 12869 16352
rect 12933 16288 12949 16352
rect 13013 16288 13021 16352
rect 12701 16282 13021 16288
rect 12701 16046 12743 16282
rect 12979 16046 13021 16282
rect 12701 15264 13021 16046
rect 12701 15200 12709 15264
rect 12773 15200 12789 15264
rect 12853 15200 12869 15264
rect 12933 15200 12949 15264
rect 13013 15200 13021 15264
rect 12701 14176 13021 15200
rect 12701 14112 12709 14176
rect 12773 14112 12789 14176
rect 12853 14112 12869 14176
rect 12933 14112 12949 14176
rect 13013 14112 13021 14176
rect 12701 13088 13021 14112
rect 12701 13024 12709 13088
rect 12773 13024 12789 13088
rect 12853 13024 12869 13088
rect 12933 13024 12949 13088
rect 13013 13024 13021 13088
rect 12701 12474 13021 13024
rect 12701 12238 12743 12474
rect 12979 12238 13021 12474
rect 12701 12000 13021 12238
rect 12701 11936 12709 12000
rect 12773 11936 12789 12000
rect 12853 11936 12869 12000
rect 12933 11936 12949 12000
rect 13013 11936 13021 12000
rect 12701 10912 13021 11936
rect 12701 10848 12709 10912
rect 12773 10848 12789 10912
rect 12853 10848 12869 10912
rect 12933 10848 12949 10912
rect 13013 10848 13021 10912
rect 12701 9824 13021 10848
rect 12701 9760 12709 9824
rect 12773 9760 12789 9824
rect 12853 9760 12869 9824
rect 12933 9760 12949 9824
rect 13013 9760 13021 9824
rect 12701 8736 13021 9760
rect 12701 8672 12709 8736
rect 12773 8672 12789 8736
rect 12853 8672 12869 8736
rect 12933 8672 12949 8736
rect 13013 8672 13021 8736
rect 12701 8666 13021 8672
rect 12701 8430 12743 8666
rect 12979 8430 13021 8666
rect 12701 7648 13021 8430
rect 12701 7584 12709 7648
rect 12773 7584 12789 7648
rect 12853 7584 12869 7648
rect 12933 7584 12949 7648
rect 13013 7584 13021 7648
rect 12701 6560 13021 7584
rect 12701 6496 12709 6560
rect 12773 6496 12789 6560
rect 12853 6496 12869 6560
rect 12933 6496 12949 6560
rect 13013 6496 13021 6560
rect 12701 5472 13021 6496
rect 12701 5408 12709 5472
rect 12773 5408 12789 5472
rect 12853 5408 12869 5472
rect 12933 5408 12949 5472
rect 13013 5408 13021 5472
rect 12701 4858 13021 5408
rect 12701 4622 12743 4858
rect 12979 4622 13021 4858
rect 12701 4384 13021 4622
rect 12701 4320 12709 4384
rect 12773 4320 12789 4384
rect 12853 4320 12869 4384
rect 12933 4320 12949 4384
rect 13013 4320 13021 4384
rect 12701 3296 13021 4320
rect 12701 3232 12709 3296
rect 12773 3232 12789 3296
rect 12853 3232 12869 3296
rect 12933 3232 12949 3296
rect 13013 3232 13021 3296
rect 12701 2208 13021 3232
rect 12701 2144 12709 2208
rect 12773 2144 12789 2208
rect 12853 2144 12869 2208
rect 12933 2144 12949 2208
rect 13013 2144 13021 2208
rect 12701 2128 13021 2144
rect 16480 16896 16800 17456
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 15622 16800 15744
rect 16480 15386 16522 15622
rect 16758 15386 16800 15622
rect 16480 14720 16800 15386
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11814 16800 12480
rect 16480 11578 16522 11814
rect 16758 11578 16800 11814
rect 16480 11456 16800 11578
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 8006 16800 8128
rect 16480 7770 16522 8006
rect 16758 7770 16800 8006
rect 16480 7104 16800 7770
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 4198 16800 4864
rect 16480 3962 16522 4198
rect 16758 3962 16800 4198
rect 16480 3840 16800 3962
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 17140 17440 17460 17456
rect 17140 17376 17148 17440
rect 17212 17376 17228 17440
rect 17292 17376 17308 17440
rect 17372 17376 17388 17440
rect 17452 17376 17460 17440
rect 17140 16352 17460 17376
rect 17140 16288 17148 16352
rect 17212 16288 17228 16352
rect 17292 16288 17308 16352
rect 17372 16288 17388 16352
rect 17452 16288 17460 16352
rect 17140 16282 17460 16288
rect 17140 16046 17182 16282
rect 17418 16046 17460 16282
rect 17140 15264 17460 16046
rect 17140 15200 17148 15264
rect 17212 15200 17228 15264
rect 17292 15200 17308 15264
rect 17372 15200 17388 15264
rect 17452 15200 17460 15264
rect 17140 14176 17460 15200
rect 17140 14112 17148 14176
rect 17212 14112 17228 14176
rect 17292 14112 17308 14176
rect 17372 14112 17388 14176
rect 17452 14112 17460 14176
rect 17140 13088 17460 14112
rect 17140 13024 17148 13088
rect 17212 13024 17228 13088
rect 17292 13024 17308 13088
rect 17372 13024 17388 13088
rect 17452 13024 17460 13088
rect 17140 12474 17460 13024
rect 17140 12238 17182 12474
rect 17418 12238 17460 12474
rect 17140 12000 17460 12238
rect 17140 11936 17148 12000
rect 17212 11936 17228 12000
rect 17292 11936 17308 12000
rect 17372 11936 17388 12000
rect 17452 11936 17460 12000
rect 17140 10912 17460 11936
rect 17140 10848 17148 10912
rect 17212 10848 17228 10912
rect 17292 10848 17308 10912
rect 17372 10848 17388 10912
rect 17452 10848 17460 10912
rect 17140 9824 17460 10848
rect 17140 9760 17148 9824
rect 17212 9760 17228 9824
rect 17292 9760 17308 9824
rect 17372 9760 17388 9824
rect 17452 9760 17460 9824
rect 17140 8736 17460 9760
rect 17140 8672 17148 8736
rect 17212 8672 17228 8736
rect 17292 8672 17308 8736
rect 17372 8672 17388 8736
rect 17452 8672 17460 8736
rect 17140 8666 17460 8672
rect 17140 8430 17182 8666
rect 17418 8430 17460 8666
rect 17140 7648 17460 8430
rect 17140 7584 17148 7648
rect 17212 7584 17228 7648
rect 17292 7584 17308 7648
rect 17372 7584 17388 7648
rect 17452 7584 17460 7648
rect 17140 6560 17460 7584
rect 17140 6496 17148 6560
rect 17212 6496 17228 6560
rect 17292 6496 17308 6560
rect 17372 6496 17388 6560
rect 17452 6496 17460 6560
rect 17140 5472 17460 6496
rect 17140 5408 17148 5472
rect 17212 5408 17228 5472
rect 17292 5408 17308 5472
rect 17372 5408 17388 5472
rect 17452 5408 17460 5472
rect 17140 4858 17460 5408
rect 17140 4622 17182 4858
rect 17418 4622 17460 4858
rect 17140 4384 17460 4622
rect 17140 4320 17148 4384
rect 17212 4320 17228 4384
rect 17292 4320 17308 4384
rect 17372 4320 17388 4384
rect 17452 4320 17460 4384
rect 17140 3296 17460 4320
rect 17140 3232 17148 3296
rect 17212 3232 17228 3296
rect 17292 3232 17308 3296
rect 17372 3232 17388 3296
rect 17452 3232 17460 3296
rect 17140 2208 17460 3232
rect 17140 2144 17148 2208
rect 17212 2144 17228 2208
rect 17292 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17460 2208
rect 17140 2128 17460 2144
<< via4 >>
rect 3205 15386 3441 15622
rect 3205 11578 3441 11814
rect 3205 7770 3441 8006
rect 3205 3962 3441 4198
rect 3865 16046 4101 16282
rect 3865 12238 4101 12474
rect 3865 8430 4101 8666
rect 3865 4622 4101 4858
rect 7644 15386 7880 15622
rect 7644 11578 7880 11814
rect 7644 7770 7880 8006
rect 7644 3962 7880 4198
rect 8304 16046 8540 16282
rect 8304 12238 8540 12474
rect 8304 8430 8540 8666
rect 8304 4622 8540 4858
rect 12083 15386 12319 15622
rect 12083 11578 12319 11814
rect 12083 7770 12319 8006
rect 12083 3962 12319 4198
rect 12743 16046 12979 16282
rect 12743 12238 12979 12474
rect 12743 8430 12979 8666
rect 12743 4622 12979 4858
rect 16522 15386 16758 15622
rect 16522 11578 16758 11814
rect 16522 7770 16758 8006
rect 16522 3962 16758 4198
rect 17182 16046 17418 16282
rect 17182 12238 17418 12474
rect 17182 8430 17418 8666
rect 17182 4622 17418 4858
<< metal5 >>
rect 1056 16282 18908 16324
rect 1056 16046 3865 16282
rect 4101 16046 8304 16282
rect 8540 16046 12743 16282
rect 12979 16046 17182 16282
rect 17418 16046 18908 16282
rect 1056 16004 18908 16046
rect 1056 15622 18908 15664
rect 1056 15386 3205 15622
rect 3441 15386 7644 15622
rect 7880 15386 12083 15622
rect 12319 15386 16522 15622
rect 16758 15386 18908 15622
rect 1056 15344 18908 15386
rect 1056 12474 18908 12516
rect 1056 12238 3865 12474
rect 4101 12238 8304 12474
rect 8540 12238 12743 12474
rect 12979 12238 17182 12474
rect 17418 12238 18908 12474
rect 1056 12196 18908 12238
rect 1056 11814 18908 11856
rect 1056 11578 3205 11814
rect 3441 11578 7644 11814
rect 7880 11578 12083 11814
rect 12319 11578 16522 11814
rect 16758 11578 18908 11814
rect 1056 11536 18908 11578
rect 1056 8666 18908 8708
rect 1056 8430 3865 8666
rect 4101 8430 8304 8666
rect 8540 8430 12743 8666
rect 12979 8430 17182 8666
rect 17418 8430 18908 8666
rect 1056 8388 18908 8430
rect 1056 8006 18908 8048
rect 1056 7770 3205 8006
rect 3441 7770 7644 8006
rect 7880 7770 12083 8006
rect 12319 7770 16522 8006
rect 16758 7770 18908 8006
rect 1056 7728 18908 7770
rect 1056 4858 18908 4900
rect 1056 4622 3865 4858
rect 4101 4622 8304 4858
rect 8540 4622 12743 4858
rect 12979 4622 17182 4858
rect 17418 4622 18908 4858
rect 1056 4580 18908 4622
rect 1056 4198 18908 4240
rect 1056 3962 3205 4198
rect 3441 3962 7644 4198
rect 7880 3962 12083 4198
rect 12319 3962 16522 4198
rect 16758 3962 18908 4198
rect 1056 3920 18908 3962
use sky130_fd_sc_hd__nor2_1  _10_
timestamp 0
transform 1 0 18216 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _11_
timestamp 0
transform -1 0 8188 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _12_
timestamp 0
transform -1 0 18492 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _13_
timestamp 0
transform 1 0 5520 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _14_
timestamp 0
transform -1 0 9476 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _16_
timestamp 0
transform -1 0 14260 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _17_
timestamp 0
transform -1 0 15824 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 0
transform 1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _19_
timestamp 0
transform -1 0 18032 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_2  _20_
timestamp 0
transform -1 0 15364 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _21_
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 0
transform 1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _24_
timestamp 0
transform -1 0 4048 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _25_
timestamp 0
transform 1 0 3864 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 0
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 0
transform 1 0 3956 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 0
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_189
timestamp 0
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 0
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_189
timestamp 0
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_35
timestamp 0
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_59
timestamp 0
transform 1 0 6532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_71
timestamp 0
transform 1 0 7636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_7
timestamp 0
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_19
timestamp 0
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_31
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_43
timestamp 0
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 0
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_7
timestamp 0
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_19
timestamp 0
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_170
timestamp 0
transform 1 0 16744 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_182
timestamp 0
transform 1 0 17848 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_7
timestamp 0
transform 1 0 1748 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_19
timestamp 0
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_31
timestamp 0
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_189
timestamp 0
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_189
timestamp 0
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_7
timestamp 0
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_19
timestamp 0
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_31
timestamp 0
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_43
timestamp 0
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_77
timestamp 0
transform 1 0 8188 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_89
timestamp 0
transform 1 0 9292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_101
timestamp 0
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 0
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_143
timestamp 0
transform 1 0 14260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_155
timestamp 0
transform 1 0 15364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 0
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_7
timestamp 0
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_19
timestamp 0
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_80
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_91
timestamp 0
transform 1 0 9476 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_103
timestamp 0
transform 1 0 10580 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_115
timestamp 0
transform 1 0 11684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_127
timestamp 0
transform 1 0 12788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 0
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_18
timestamp 0
transform 1 0 2760 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_24
timestamp 0
transform 1 0 3312 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_32
timestamp 0
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_44
timestamp 0
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_181
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_189
timestamp 0
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 0
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 0
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_189
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_78
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_90
timestamp 0
transform 1 0 9384 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 0
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 0
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 0
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_6
timestamp 0
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 0
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 0
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 0
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_189
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_7
timestamp 0
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_19
timestamp 0
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_31
timestamp 0
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_43
timestamp 0
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_189
timestamp 0
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_7
timestamp 0
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_19
timestamp 0
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_189
timestamp 0
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_7
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_19
timestamp 0
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_31
timestamp 0
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 0
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 0
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 0
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 0
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_7
timestamp 0
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_19
timestamp 0
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_31
timestamp 0
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_43
timestamp 0
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_189
timestamp 0
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_7
timestamp 0
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 0
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_47
timestamp 0
transform 1 0 5428 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_57
timestamp 0
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_69
timestamp 0
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 0
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_189
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_7
timestamp 0
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_19
timestamp 0
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_31
timestamp 0
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_43
timestamp 0
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_87
timestamp 0
transform 1 0 9108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_99
timestamp 0
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_185
timestamp 0
transform 1 0 18124 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 0
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_7
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_19
timestamp 0
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_181
timestamp 0
transform 1 0 17756 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 0
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_7
timestamp 0
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_19
timestamp 0
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_160
timestamp 0
transform 1 0 15824 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_172
timestamp 0
transform 1 0 16928 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_184
timestamp 0
transform 1 0 18032 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_184
timestamp 0
transform 1 0 18032 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_34
timestamp 0
transform 1 0 4232 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_46
timestamp 0
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_58
timestamp 0
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_70
timestamp 0
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_82
timestamp 0
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_147
timestamp 0
transform 1 0 14628 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_155
timestamp 0
transform 1 0 15364 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_167
timestamp 0
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_179
timestamp 0
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_187
timestamp 0
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 0
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 0
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 0
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_63
timestamp 0
transform 1 0 6900 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_75
timestamp 0
transform 1 0 8004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_83
timestamp 0
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_85
timestamp 0
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_97
timestamp 0
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 0
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 0
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 0
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 0
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 0
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 0
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 0
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 0
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 0
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 0
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 0
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 0
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 0
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 0
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 0
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 0
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 0
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
rlabel metal1 s 9982 17408 9982 17408 4 VGND
rlabel metal1 s 9982 16864 9982 16864 4 VPWR
rlabel metal1 s 17112 5678 17112 5678 4 _00_
rlabel metal2 s 18446 11016 18446 11016 4 _01_
rlabel metal1 s 6440 17034 6440 17034 4 _02_
rlabel metal1 s 8418 7888 8418 7888 4 _03_
rlabel metal2 s 17066 11628 17066 11628 4 _04_
rlabel metal1 s 5842 2380 5842 2380 4 _05_
rlabel metal1 s 9476 9486 9476 9486 4 _06_
rlabel metal1 s 7452 17306 7452 17306 4 _07_
rlabel metal1 s 8648 9622 8648 9622 4 _08_
rlabel metal2 s 13846 5066 13846 5066 4 _09_
rlabel metal1 s 4968 4590 4968 4590 4 net1
rlabel metal1 s 1794 14382 1794 14382 4 net10
rlabel metal2 s 3726 9622 3726 9622 4 net11
rlabel metal1 s 4324 5678 4324 5678 4 net12
rlabel metal1 s 3772 2618 3772 2618 4 net13
rlabel metal1 s 1748 6290 1748 6290 4 net14
rlabel metal1 s 4301 13906 4301 13906 4 net15
rlabel metal1 s 2254 7854 2254 7854 4 net16
rlabel metal1 s 3818 4658 3818 4658 4 net2
rlabel metal2 s 5731 13294 5731 13294 4 net3
rlabel metal1 s 5198 13226 5198 13226 4 net4
rlabel metal1 s 6394 17204 6394 17204 4 net5
rlabel metal1 s 5957 16966 5957 16966 4 net6
rlabel metal1 s 4232 9146 4232 9146 4 net7
rlabel metal1 s 2714 8466 2714 8466 4 net8
rlabel metal1 s 3818 16422 3818 16422 4 net9
rlabel metal3 s 0 4768 800 4888 4 x[0]
port 3 nsew
rlabel metal3 s 0 10208 800 10328 4 x[1]
port 4 nsew
rlabel metal3 s 1096 10948 1096 10948 4 x[2]
rlabel metal3 s 1050 9588 1050 9588 4 x[3]
rlabel metal3 s 1096 6868 1096 6868 4 x[4]
rlabel metal3 s 1096 12308 1096 12308 4 x[5]
rlabel metal3 s 0 8848 800 8968 4 x[6]
port 9 nsew
rlabel metal3 s 1050 8228 1050 8228 4 x[7]
rlabel metal3 s 0 12928 800 13048 4 y[0]
port 11 nsew
rlabel metal3 s 0 14288 800 14408 4 y[1]
port 12 nsew
rlabel metal3 s 0 11568 800 11688 4 y[2]
port 13 nsew
rlabel metal3 s 1096 5508 1096 5508 4 y[3]
rlabel metal3 s 1096 15028 1096 15028 4 y[4]
rlabel metal3 s 0 6128 800 6248 4 y[5]
port 16 nsew
rlabel metal3 s 1096 13668 1096 13668 4 y[6]
rlabel metal3 s 0 7488 800 7608 4 y[7]
port 18 nsew
flabel metal5 s 1056 16004 18908 16324 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 12196 18908 12516 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8388 18908 8708 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 4580 18908 4900 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 17140 2128 17460 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12701 2128 13021 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8262 2128 8582 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3823 2128 4143 17456 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 15344 18908 15664 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 11536 18908 11856 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 7728 18908 8048 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3920 18908 4240 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 16480 2128 16800 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12041 2128 12361 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7602 2128 7922 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3163 2128 3483 17456 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 400 4828 400 4828 0 FreeSans 600 0 0 0 x[0]
flabel metal3 s 400 10268 400 10268 0 FreeSans 600 0 0 0 x[1]
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 x[2]
port 5 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 x[3]
port 6 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 x[4]
port 7 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 x[5]
port 8 nsew
flabel metal3 s 400 8908 400 8908 0 FreeSans 600 0 0 0 x[6]
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 x[7]
port 10 nsew
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 y[0]
flabel metal3 s 400 14348 400 14348 0 FreeSans 600 0 0 0 y[1]
flabel metal3 s 400 11628 400 11628 0 FreeSans 600 0 0 0 y[2]
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 y[3]
port 14 nsew
flabel metal3 s 0 14968 800 15088 0 FreeSans 600 0 0 0 y[4]
port 15 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 y[5]
flabel metal3 s 0 13608 800 13728 0 FreeSans 600 0 0 0 y[6]
port 17 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 y[7]
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
